// Benchmark "top" written by ABC on Wed Jan 17 21:32:50 2024

module top ( 
    i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_, i_10_,
    i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_,
    i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_, i_24_,
    i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_, i_32_,
    i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_, i_19_,
    i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_, i_38_,
    i_29_, i_51_, i_44_, i_37_,
    o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_  );
  input  i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_,
    i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_,
    i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_,
    i_24_, i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_,
    i_32_, i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_,
    i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_,
    i_38_, i_29_, i_51_, i_44_, i_37_;
  output o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_;
  wire new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1156_, new_n1157_, new_n1158_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1170_, new_n1171_, new_n1172_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1236_, new_n1237_, new_n1238_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1246_, new_n1247_, new_n1248_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1270_,
    new_n1271_, new_n1272_, new_n1274_, new_n1275_, new_n1276_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1296_;
  nor2 g0000(.a(i_24_), .b(i_25_), .O(new_n131_));
  inv1 g0001(.a(new_n131_), .O(new_n132_));
  nor2 g0002(.a(new_n132_), .b(i_26_), .O(new_n133_));
  inv1 g0003(.a(new_n133_), .O(new_n134_));
  inv1 g0004(.a(i_29_), .O(new_n135_));
  nor2 g0005(.a(new_n135_), .b(i_28_), .O(new_n136_));
  inv1 g0006(.a(new_n136_), .O(new_n137_));
  nor2 g0007(.a(new_n135_), .b(i_30_), .O(new_n138_));
  inv1 g0008(.a(new_n138_), .O(new_n139_));
  nor2 g0009(.a(new_n139_), .b(new_n137_), .O(new_n140_));
  inv1 g0010(.a(new_n140_), .O(new_n141_));
  nor2 g0011(.a(new_n141_), .b(new_n134_), .O(new_n142_));
  inv1 g0012(.a(new_n142_), .O(new_n143_));
  nor2 g0013(.a(i_33_), .b(i_34_), .O(new_n144_));
  inv1 g0014(.a(new_n144_), .O(new_n145_));
  nor2 g0015(.a(new_n145_), .b(i_31_), .O(new_n146_));
  inv1 g0016(.a(new_n146_), .O(new_n147_));
  nor2 g0017(.a(new_n147_), .b(new_n143_), .O(new_n148_));
  inv1 g0018(.a(new_n148_), .O(new_n149_));
  nor2 g0019(.a(i_22_), .b(i_18_), .O(new_n150_));
  inv1 g0020(.a(new_n150_), .O(new_n151_));
  nor2 g0021(.a(new_n151_), .b(i_17_), .O(new_n152_));
  inv1 g0022(.a(new_n152_), .O(new_n153_));
  nor2 g0023(.a(i_37_), .b(i_39_), .O(new_n154_));
  inv1 g0024(.a(new_n154_), .O(new_n155_));
  nor2 g0025(.a(new_n155_), .b(i_35_), .O(new_n156_));
  inv1 g0026(.a(new_n156_), .O(new_n157_));
  nor2 g0027(.a(new_n157_), .b(new_n153_), .O(new_n158_));
  inv1 g0028(.a(new_n158_), .O(new_n159_));
  nor2 g0029(.a(i_15_), .b(i_14_), .O(new_n160_));
  inv1 g0030(.a(new_n160_), .O(new_n161_));
  nor2 g0031(.a(new_n161_), .b(i_11_), .O(new_n162_));
  inv1 g0032(.a(new_n162_), .O(new_n163_));
  nor2 g0033(.a(new_n163_), .b(new_n159_), .O(new_n164_));
  inv1 g0034(.a(new_n164_), .O(new_n165_));
  nor2 g0035(.a(new_n165_), .b(new_n149_), .O(new_n166_));
  inv1 g0036(.a(new_n166_), .O(new_n167_));
  nor2 g0037(.a(i_41_), .b(i_40_), .O(new_n168_));
  inv1 g0038(.a(new_n168_), .O(new_n169_));
  nor2 g0039(.a(new_n169_), .b(i_42_), .O(new_n170_));
  inv1 g0040(.a(new_n170_), .O(new_n171_));
  nor2 g0041(.a(i_47_), .b(i_46_), .O(new_n172_));
  inv1 g0042(.a(new_n172_), .O(new_n173_));
  nor2 g0043(.a(new_n173_), .b(i_43_), .O(new_n174_));
  inv1 g0044(.a(new_n174_), .O(new_n175_));
  inv1 g0045(.a(i_5_), .O(new_n176_));
  nor2 g0046(.a(i_6_), .b(i_7_), .O(new_n177_));
  inv1 g0047(.a(new_n177_), .O(new_n178_));
  nor2 g0048(.a(new_n178_), .b(new_n176_), .O(new_n179_));
  inv1 g0049(.a(new_n179_), .O(new_n180_));
  nor2 g0050(.a(new_n180_), .b(new_n175_), .O(new_n181_));
  inv1 g0051(.a(new_n181_), .O(new_n182_));
  nor2 g0052(.a(new_n182_), .b(new_n171_), .O(new_n183_));
  inv1 g0053(.a(new_n183_), .O(new_n184_));
  nor2 g0054(.a(i_55_), .b(i_56_), .O(new_n185_));
  inv1 g0055(.a(new_n185_), .O(new_n186_));
  nor2 g0056(.a(new_n186_), .b(i_54_), .O(new_n187_));
  inv1 g0057(.a(new_n187_), .O(new_n188_));
  nor2 g0058(.a(i_51_), .b(i_50_), .O(new_n189_));
  inv1 g0059(.a(new_n189_), .O(new_n190_));
  nor2 g0060(.a(new_n190_), .b(i_53_), .O(new_n191_));
  inv1 g0061(.a(new_n191_), .O(new_n192_));
  nor2 g0062(.a(new_n192_), .b(new_n188_), .O(new_n193_));
  inv1 g0063(.a(new_n193_), .O(new_n194_));
  nor2 g0064(.a(i_4_), .b(i_3_), .O(new_n195_));
  inv1 g0065(.a(new_n195_), .O(new_n196_));
  nor2 g0066(.a(new_n196_), .b(i_0_), .O(new_n197_));
  inv1 g0067(.a(new_n197_), .O(new_n198_));
  nor2 g0068(.a(i_8_), .b(i_10_), .O(new_n199_));
  inv1 g0069(.a(new_n199_), .O(new_n200_));
  nor2 g0070(.a(new_n200_), .b(i_9_), .O(new_n201_));
  inv1 g0071(.a(new_n201_), .O(new_n202_));
  nor2 g0072(.a(new_n202_), .b(new_n198_), .O(new_n203_));
  inv1 g0073(.a(new_n203_), .O(new_n204_));
  nor2 g0074(.a(i_58_), .b(i_59_), .O(new_n205_));
  inv1 g0075(.a(new_n205_), .O(new_n206_));
  nor2 g0076(.a(i_62_), .b(i_61_), .O(new_n207_));
  inv1 g0077(.a(new_n207_), .O(new_n208_));
  nor2 g0078(.a(new_n208_), .b(i_60_), .O(new_n209_));
  inv1 g0079(.a(new_n209_), .O(new_n210_));
  nor2 g0080(.a(new_n210_), .b(new_n206_), .O(new_n211_));
  inv1 g0081(.a(new_n211_), .O(new_n212_));
  nor2 g0082(.a(new_n212_), .b(new_n204_), .O(new_n213_));
  inv1 g0083(.a(new_n213_), .O(new_n214_));
  nor2 g0084(.a(new_n214_), .b(new_n194_), .O(new_n215_));
  inv1 g0085(.a(new_n215_), .O(new_n216_));
  nor2 g0086(.a(new_n216_), .b(new_n184_), .O(new_n217_));
  inv1 g0087(.a(new_n217_), .O(new_n218_));
  nor2 g0088(.a(new_n218_), .b(new_n167_), .O(o_1_));
  nor2 g0089(.a(i_8_), .b(i_7_), .O(new_n220_));
  inv1 g0090(.a(new_n220_), .O(new_n221_));
  nor2 g0091(.a(i_6_), .b(i_5_), .O(new_n222_));
  inv1 g0092(.a(new_n222_), .O(new_n223_));
  nor2 g0093(.a(new_n223_), .b(new_n196_), .O(new_n224_));
  inv1 g0094(.a(new_n224_), .O(new_n225_));
  nor2 g0095(.a(new_n225_), .b(new_n221_), .O(new_n226_));
  inv1 g0096(.a(new_n226_), .O(new_n227_));
  nor2 g0097(.a(i_2_), .b(i_1_), .O(new_n228_));
  inv1 g0098(.a(new_n228_), .O(new_n229_));
  nor2 g0099(.a(new_n229_), .b(i_0_), .O(new_n230_));
  inv1 g0100(.a(new_n230_), .O(new_n231_));
  nor2 g0101(.a(new_n231_), .b(new_n227_), .O(new_n232_));
  inv1 g0102(.a(new_n232_), .O(new_n233_));
  nor2 g0103(.a(i_25_), .b(i_28_), .O(new_n234_));
  inv1 g0104(.a(new_n234_), .O(new_n235_));
  nor2 g0105(.a(new_n235_), .b(i_24_), .O(new_n236_));
  inv1 g0106(.a(new_n236_), .O(new_n237_));
  nor2 g0107(.a(new_n151_), .b(i_26_), .O(new_n238_));
  inv1 g0108(.a(new_n238_), .O(new_n239_));
  nor2 g0109(.a(new_n239_), .b(new_n237_), .O(new_n240_));
  inv1 g0110(.a(new_n240_), .O(new_n241_));
  nor2 g0111(.a(new_n161_), .b(i_17_), .O(new_n242_));
  inv1 g0112(.a(new_n242_), .O(new_n243_));
  nor2 g0113(.a(new_n243_), .b(new_n241_), .O(new_n244_));
  inv1 g0114(.a(new_n244_), .O(new_n245_));
  nor2 g0115(.a(i_11_), .b(i_10_), .O(new_n246_));
  inv1 g0116(.a(new_n246_), .O(new_n247_));
  nor2 g0117(.a(new_n247_), .b(i_9_), .O(new_n248_));
  inv1 g0118(.a(new_n248_), .O(new_n249_));
  nor2 g0119(.a(i_31_), .b(i_30_), .O(new_n250_));
  inv1 g0120(.a(new_n250_), .O(new_n251_));
  nor2 g0121(.a(new_n251_), .b(new_n135_), .O(new_n252_));
  inv1 g0122(.a(new_n252_), .O(new_n253_));
  nor2 g0123(.a(new_n145_), .b(i_35_), .O(new_n254_));
  inv1 g0124(.a(new_n254_), .O(new_n255_));
  nor2 g0125(.a(new_n255_), .b(new_n253_), .O(new_n256_));
  inv1 g0126(.a(new_n256_), .O(new_n257_));
  nor2 g0127(.a(new_n257_), .b(new_n249_), .O(new_n258_));
  inv1 g0128(.a(new_n258_), .O(new_n259_));
  nor2 g0129(.a(new_n259_), .b(new_n245_), .O(new_n260_));
  inv1 g0130(.a(new_n260_), .O(new_n261_));
  nor2 g0131(.a(new_n261_), .b(new_n233_), .O(new_n262_));
  inv1 g0132(.a(new_n262_), .O(new_n263_));
  nor2 g0133(.a(new_n173_), .b(i_45_), .O(new_n264_));
  inv1 g0134(.a(new_n264_), .O(new_n265_));
  nor2 g0135(.a(i_39_), .b(i_40_), .O(new_n266_));
  inv1 g0136(.a(new_n266_), .O(new_n267_));
  nor2 g0137(.a(new_n267_), .b(i_41_), .O(new_n268_));
  inv1 g0138(.a(new_n268_), .O(new_n269_));
  nor2 g0139(.a(i_43_), .b(i_42_), .O(new_n270_));
  inv1 g0140(.a(new_n270_), .O(new_n271_));
  nor2 g0141(.a(new_n271_), .b(i_37_), .O(new_n272_));
  inv1 g0142(.a(new_n272_), .O(new_n273_));
  nor2 g0143(.a(new_n273_), .b(new_n269_), .O(new_n274_));
  inv1 g0144(.a(new_n274_), .O(new_n275_));
  nor2 g0145(.a(new_n275_), .b(new_n265_), .O(new_n276_));
  inv1 g0146(.a(new_n276_), .O(new_n277_));
  nor2 g0147(.a(new_n277_), .b(new_n212_), .O(new_n278_));
  inv1 g0148(.a(new_n278_), .O(new_n279_));
  inv1 g0149(.a(i_64_), .O(new_n280_));
  nor2 g0150(.a(i_49_), .b(i_50_), .O(new_n281_));
  inv1 g0151(.a(new_n281_), .O(new_n282_));
  nor2 g0152(.a(new_n282_), .b(i_48_), .O(new_n283_));
  inv1 g0153(.a(new_n283_), .O(new_n284_));
  nor2 g0154(.a(i_53_), .b(i_54_), .O(new_n285_));
  inv1 g0155(.a(new_n285_), .O(new_n286_));
  nor2 g0156(.a(new_n286_), .b(i_51_), .O(new_n287_));
  inv1 g0157(.a(new_n287_), .O(new_n288_));
  nor2 g0158(.a(new_n288_), .b(new_n284_), .O(new_n289_));
  inv1 g0159(.a(new_n289_), .O(new_n290_));
  nor2 g0160(.a(new_n186_), .b(i_57_), .O(new_n291_));
  inv1 g0161(.a(new_n291_), .O(new_n292_));
  nor2 g0162(.a(new_n292_), .b(new_n290_), .O(new_n293_));
  inv1 g0163(.a(new_n293_), .O(new_n294_));
  nor2 g0164(.a(new_n294_), .b(new_n280_), .O(new_n295_));
  inv1 g0165(.a(new_n295_), .O(new_n296_));
  nor2 g0166(.a(new_n296_), .b(new_n279_), .O(new_n297_));
  inv1 g0167(.a(new_n297_), .O(new_n298_));
  nor2 g0168(.a(new_n298_), .b(new_n263_), .O(o_19_));
  nor2 g0169(.a(i_16_), .b(i_17_), .O(new_n300_));
  inv1 g0170(.a(new_n300_), .O(new_n301_));
  nor2 g0171(.a(new_n301_), .b(i_15_), .O(new_n302_));
  inv1 g0172(.a(new_n302_), .O(new_n303_));
  nor2 g0173(.a(new_n303_), .b(new_n249_), .O(new_n304_));
  inv1 g0174(.a(new_n304_), .O(new_n305_));
  nor2 g0175(.a(i_12_), .b(i_14_), .O(new_n306_));
  inv1 g0176(.a(new_n306_), .O(new_n307_));
  nor2 g0177(.a(new_n307_), .b(i_13_), .O(new_n308_));
  inv1 g0178(.a(new_n308_), .O(new_n309_));
  nor2 g0179(.a(new_n309_), .b(new_n305_), .O(new_n310_));
  inv1 g0180(.a(new_n310_), .O(new_n311_));
  nor2 g0181(.a(new_n311_), .b(new_n233_), .O(new_n312_));
  inv1 g0182(.a(new_n312_), .O(new_n313_));
  inv1 g0183(.a(i_23_), .O(new_n314_));
  nor2 g0184(.a(i_21_), .b(new_n314_), .O(new_n315_));
  inv1 g0185(.a(new_n315_), .O(new_n316_));
  nor2 g0186(.a(new_n316_), .b(i_22_), .O(new_n317_));
  inv1 g0187(.a(new_n317_), .O(new_n318_));
  nor2 g0188(.a(new_n318_), .b(new_n134_), .O(new_n319_));
  nor2 g0189(.a(i_18_), .b(i_20_), .O(new_n320_));
  inv1 g0190(.a(new_n320_), .O(new_n321_));
  nor2 g0191(.a(new_n321_), .b(i_19_), .O(new_n322_));
  inv1 g0192(.a(new_n322_), .O(new_n323_));
  nor2 g0193(.a(i_21_), .b(i_24_), .O(new_n324_));
  inv1 g0194(.a(new_n324_), .O(new_n325_));
  nor2 g0195(.a(new_n325_), .b(i_22_), .O(new_n326_));
  inv1 g0196(.a(new_n326_), .O(new_n327_));
  nor2 g0197(.a(new_n327_), .b(new_n134_), .O(new_n328_));
  inv1 g0198(.a(new_n328_), .O(new_n329_));
  nor2 g0199(.a(new_n329_), .b(new_n323_), .O(new_n330_));
  inv1 g0200(.a(new_n330_), .O(new_n331_));
  nor2 g0201(.a(new_n331_), .b(new_n319_), .O(new_n332_));
  inv1 g0202(.a(new_n332_), .O(new_n333_));
  nor2 g0203(.a(new_n333_), .b(new_n313_), .O(new_n334_));
  inv1 g0204(.a(new_n334_), .O(new_n335_));
  inv1 g0205(.a(i_27_), .O(new_n336_));
  nor2 g0206(.a(i_32_), .b(new_n336_), .O(new_n337_));
  inv1 g0207(.a(new_n337_), .O(new_n338_));
  nor2 g0208(.a(i_44_), .b(i_38_), .O(new_n339_));
  inv1 g0209(.a(new_n339_), .O(new_n340_));
  nor2 g0210(.a(new_n340_), .b(new_n338_), .O(new_n341_));
  inv1 g0211(.a(new_n341_), .O(new_n342_));
  nor2 g0212(.a(i_64_), .b(i_63_), .O(new_n343_));
  inv1 g0213(.a(new_n343_), .O(new_n344_));
  nor2 g0214(.a(i_36_), .b(i_31_), .O(new_n345_));
  inv1 g0215(.a(new_n345_), .O(new_n346_));
  nor2 g0216(.a(new_n346_), .b(new_n344_), .O(new_n347_));
  inv1 g0217(.a(new_n347_), .O(new_n348_));
  nor2 g0218(.a(new_n348_), .b(new_n342_), .O(new_n349_));
  inv1 g0219(.a(new_n349_), .O(new_n350_));
  nor2 g0220(.a(new_n350_), .b(new_n275_), .O(new_n351_));
  inv1 g0221(.a(new_n351_), .O(new_n352_));
  nor2 g0222(.a(new_n284_), .b(new_n265_), .O(new_n353_));
  inv1 g0223(.a(new_n353_), .O(new_n354_));
  nor2 g0224(.a(new_n255_), .b(new_n141_), .O(new_n355_));
  inv1 g0225(.a(new_n355_), .O(new_n356_));
  nor2 g0226(.a(new_n356_), .b(new_n354_), .O(new_n357_));
  inv1 g0227(.a(new_n357_), .O(new_n358_));
  nor2 g0228(.a(new_n206_), .b(i_57_), .O(new_n359_));
  inv1 g0229(.a(new_n359_), .O(new_n360_));
  nor2 g0230(.a(new_n360_), .b(new_n210_), .O(new_n361_));
  inv1 g0231(.a(new_n361_), .O(new_n362_));
  nor2 g0232(.a(i_52_), .b(i_53_), .O(new_n363_));
  inv1 g0233(.a(new_n363_), .O(new_n364_));
  nor2 g0234(.a(new_n364_), .b(i_51_), .O(new_n365_));
  inv1 g0235(.a(new_n365_), .O(new_n366_));
  nor2 g0236(.a(new_n366_), .b(new_n188_), .O(new_n367_));
  inv1 g0237(.a(new_n367_), .O(new_n368_));
  nor2 g0238(.a(new_n368_), .b(new_n362_), .O(new_n369_));
  inv1 g0239(.a(new_n369_), .O(new_n370_));
  nor2 g0240(.a(new_n370_), .b(new_n358_), .O(new_n371_));
  inv1 g0241(.a(new_n371_), .O(new_n372_));
  nor2 g0242(.a(new_n372_), .b(new_n352_), .O(new_n373_));
  inv1 g0243(.a(new_n373_), .O(new_n374_));
  nor2 g0244(.a(new_n374_), .b(new_n335_), .O(o_2_));
  nor2 g0245(.a(i_56_), .b(i_58_), .O(new_n376_));
  inv1 g0246(.a(new_n376_), .O(new_n377_));
  nor2 g0247(.a(new_n210_), .b(i_59_), .O(new_n378_));
  inv1 g0248(.a(new_n378_), .O(new_n379_));
  nor2 g0249(.a(new_n379_), .b(new_n377_), .O(new_n380_));
  inv1 g0250(.a(new_n380_), .O(new_n381_));
  nor2 g0251(.a(new_n190_), .b(i_47_), .O(new_n382_));
  inv1 g0252(.a(new_n382_), .O(new_n383_));
  nor2 g0253(.a(i_54_), .b(i_55_), .O(new_n384_));
  inv1 g0254(.a(new_n384_), .O(new_n385_));
  nor2 g0255(.a(new_n385_), .b(i_53_), .O(new_n386_));
  inv1 g0256(.a(new_n386_), .O(new_n387_));
  nor2 g0257(.a(new_n387_), .b(new_n171_), .O(new_n388_));
  inv1 g0258(.a(new_n388_), .O(new_n389_));
  nor2 g0259(.a(new_n389_), .b(new_n383_), .O(new_n390_));
  inv1 g0260(.a(new_n390_), .O(new_n391_));
  nor2 g0261(.a(i_43_), .b(i_46_), .O(new_n392_));
  inv1 g0262(.a(new_n392_), .O(new_n393_));
  inv1 g0263(.a(i_45_), .O(new_n394_));
  nor2 g0264(.a(new_n394_), .b(i_5_), .O(new_n395_));
  inv1 g0265(.a(new_n395_), .O(new_n396_));
  nor2 g0266(.a(new_n396_), .b(new_n178_), .O(new_n397_));
  inv1 g0267(.a(new_n397_), .O(new_n398_));
  nor2 g0268(.a(new_n398_), .b(new_n393_), .O(new_n399_));
  inv1 g0269(.a(new_n399_), .O(new_n400_));
  nor2 g0270(.a(new_n400_), .b(new_n204_), .O(new_n401_));
  inv1 g0271(.a(new_n401_), .O(new_n402_));
  nor2 g0272(.a(new_n402_), .b(new_n391_), .O(new_n403_));
  inv1 g0273(.a(new_n403_), .O(new_n404_));
  nor2 g0274(.a(new_n404_), .b(new_n381_), .O(new_n405_));
  inv1 g0275(.a(new_n405_), .O(new_n406_));
  nor2 g0276(.a(new_n406_), .b(new_n167_), .O(o_0_));
  nor2 g0277(.a(new_n161_), .b(i_10_), .O(new_n408_));
  inv1 g0278(.a(new_n408_), .O(new_n409_));
  nor2 g0279(.a(new_n137_), .b(i_37_), .O(new_n410_));
  inv1 g0280(.a(new_n410_), .O(new_n411_));
  nor2 g0281(.a(new_n411_), .b(i_43_), .O(new_n412_));
  inv1 g0282(.a(new_n412_), .O(new_n413_));
  nor2 g0283(.a(new_n413_), .b(new_n267_), .O(new_n414_));
  inv1 g0284(.a(new_n414_), .O(new_n415_));
  nor2 g0285(.a(new_n415_), .b(new_n409_), .O(new_n416_));
  inv1 g0286(.a(new_n416_), .O(new_n417_));
  inv1 g0287(.a(i_60_), .O(new_n418_));
  nor2 g0288(.a(i_58_), .b(i_50_), .O(new_n419_));
  inv1 g0289(.a(new_n419_), .O(new_n420_));
  nor2 g0290(.a(new_n420_), .b(i_46_), .O(new_n421_));
  inv1 g0291(.a(new_n421_), .O(new_n422_));
  nor2 g0292(.a(new_n422_), .b(new_n418_), .O(new_n423_));
  inv1 g0293(.a(new_n423_), .O(new_n424_));
  nor2 g0294(.a(new_n424_), .b(new_n417_), .O(o_29_));
  nor2 g0295(.a(i_43_), .b(i_40_), .O(new_n426_));
  inv1 g0296(.a(new_n426_), .O(new_n427_));
  nor2 g0297(.a(new_n427_), .b(i_39_), .O(new_n428_));
  inv1 g0298(.a(new_n428_), .O(new_n429_));
  nor2 g0299(.a(new_n429_), .b(new_n163_), .O(new_n430_));
  inv1 g0300(.a(new_n430_), .O(new_n431_));
  nor2 g0301(.a(new_n139_), .b(i_37_), .O(new_n432_));
  inv1 g0302(.a(new_n432_), .O(new_n433_));
  nor2 g0303(.a(i_46_), .b(i_50_), .O(new_n434_));
  inv1 g0304(.a(new_n434_), .O(new_n435_));
  nor2 g0305(.a(new_n435_), .b(i_47_), .O(new_n436_));
  inv1 g0306(.a(new_n436_), .O(new_n437_));
  nor2 g0307(.a(new_n437_), .b(new_n237_), .O(new_n438_));
  inv1 g0308(.a(new_n438_), .O(new_n439_));
  nor2 g0309(.a(new_n439_), .b(new_n433_), .O(new_n440_));
  inv1 g0310(.a(new_n440_), .O(new_n441_));
  nor2 g0311(.a(new_n441_), .b(new_n431_), .O(new_n442_));
  inv1 g0312(.a(new_n442_), .O(new_n443_));
  nor2 g0313(.a(i_60_), .b(i_58_), .O(new_n444_));
  inv1 g0314(.a(new_n444_), .O(new_n445_));
  nor2 g0315(.a(new_n445_), .b(i_56_), .O(new_n446_));
  inv1 g0316(.a(new_n446_), .O(new_n447_));
  inv1 g0317(.a(i_7_), .O(new_n448_));
  nor2 g0318(.a(new_n200_), .b(new_n448_), .O(new_n449_));
  inv1 g0319(.a(new_n449_), .O(new_n450_));
  nor2 g0320(.a(new_n450_), .b(new_n447_), .O(new_n451_));
  inv1 g0321(.a(new_n451_), .O(new_n452_));
  nor2 g0322(.a(new_n452_), .b(new_n443_), .O(o_60_));
  nor2 g0323(.a(new_n247_), .b(i_14_), .O(new_n454_));
  inv1 g0324(.a(new_n454_), .O(new_n455_));
  nor2 g0325(.a(new_n221_), .b(i_6_), .O(new_n456_));
  inv1 g0326(.a(new_n456_), .O(new_n457_));
  nor2 g0327(.a(new_n457_), .b(new_n198_), .O(new_n458_));
  inv1 g0328(.a(new_n458_), .O(new_n459_));
  nor2 g0329(.a(new_n459_), .b(new_n455_), .O(new_n460_));
  inv1 g0330(.a(new_n460_), .O(new_n461_));
  nor2 g0331(.a(new_n151_), .b(i_15_), .O(new_n462_));
  inv1 g0332(.a(new_n462_), .O(new_n463_));
  nor2 g0333(.a(new_n463_), .b(new_n143_), .O(new_n464_));
  inv1 g0334(.a(new_n464_), .O(new_n465_));
  nor2 g0335(.a(new_n465_), .b(new_n461_), .O(new_n466_));
  inv1 g0336(.a(new_n466_), .O(new_n467_));
  nor2 g0337(.a(new_n175_), .b(new_n157_), .O(new_n468_));
  inv1 g0338(.a(new_n468_), .O(new_n469_));
  nor2 g0339(.a(new_n445_), .b(new_n186_), .O(new_n470_));
  inv1 g0340(.a(new_n470_), .O(new_n471_));
  inv1 g0341(.a(i_42_), .O(new_n472_));
  nor2 g0342(.a(new_n208_), .b(new_n472_), .O(new_n473_));
  inv1 g0343(.a(new_n473_), .O(new_n474_));
  nor2 g0344(.a(new_n190_), .b(new_n169_), .O(new_n475_));
  inv1 g0345(.a(new_n475_), .O(new_n476_));
  nor2 g0346(.a(new_n476_), .b(new_n474_), .O(new_n477_));
  inv1 g0347(.a(new_n477_), .O(new_n478_));
  nor2 g0348(.a(new_n478_), .b(new_n471_), .O(new_n479_));
  inv1 g0349(.a(new_n479_), .O(new_n480_));
  nor2 g0350(.a(new_n480_), .b(new_n469_), .O(new_n481_));
  inv1 g0351(.a(new_n481_), .O(new_n482_));
  nor2 g0352(.a(new_n482_), .b(new_n467_), .O(o_39_));
  nor2 g0353(.a(new_n190_), .b(i_55_), .O(new_n484_));
  inv1 g0354(.a(new_n484_), .O(new_n485_));
  nor2 g0355(.a(new_n485_), .b(new_n171_), .O(new_n486_));
  inv1 g0356(.a(new_n486_), .O(new_n487_));
  inv1 g0357(.a(i_59_), .O(new_n488_));
  nor2 g0358(.a(new_n377_), .b(new_n488_), .O(new_n489_));
  inv1 g0359(.a(new_n489_), .O(new_n490_));
  nor2 g0360(.a(new_n490_), .b(new_n210_), .O(new_n491_));
  inv1 g0361(.a(new_n491_), .O(new_n492_));
  nor2 g0362(.a(new_n492_), .b(new_n469_), .O(new_n493_));
  inv1 g0363(.a(new_n493_), .O(new_n494_));
  nor2 g0364(.a(new_n494_), .b(new_n487_), .O(new_n495_));
  inv1 g0365(.a(new_n495_), .O(new_n496_));
  nor2 g0366(.a(new_n496_), .b(new_n467_), .O(o_38_));
  nor2 g0367(.a(new_n445_), .b(new_n393_), .O(new_n498_));
  inv1 g0368(.a(new_n498_), .O(new_n499_));
  nor2 g0369(.a(new_n135_), .b(i_15_), .O(new_n500_));
  inv1 g0370(.a(new_n500_), .O(new_n501_));
  nor2 g0371(.a(i_14_), .b(i_10_), .O(new_n502_));
  inv1 g0372(.a(new_n502_), .O(new_n503_));
  nor2 g0373(.a(new_n503_), .b(new_n501_), .O(new_n504_));
  inv1 g0374(.a(new_n504_), .O(new_n505_));
  nor2 g0375(.a(new_n505_), .b(new_n499_), .O(new_n506_));
  inv1 g0376(.a(new_n506_), .O(new_n507_));
  inv1 g0377(.a(i_24_), .O(new_n508_));
  nor2 g0378(.a(i_40_), .b(i_50_), .O(new_n509_));
  inv1 g0379(.a(new_n509_), .O(new_n510_));
  nor2 g0380(.a(new_n510_), .b(new_n508_), .O(new_n511_));
  inv1 g0381(.a(new_n511_), .O(new_n512_));
  nor2 g0382(.a(new_n235_), .b(new_n155_), .O(new_n513_));
  inv1 g0383(.a(new_n513_), .O(new_n514_));
  nor2 g0384(.a(new_n514_), .b(new_n512_), .O(new_n515_));
  inv1 g0385(.a(new_n515_), .O(new_n516_));
  nor2 g0386(.a(new_n516_), .b(new_n507_), .O(o_25_));
  nor2 g0387(.a(new_n447_), .b(i_50_), .O(new_n518_));
  inv1 g0388(.a(new_n518_), .O(new_n519_));
  nor2 g0389(.a(new_n519_), .b(i_62_), .O(new_n520_));
  inv1 g0390(.a(new_n520_), .O(new_n521_));
  nor2 g0391(.a(new_n521_), .b(new_n175_), .O(new_n522_));
  inv1 g0392(.a(new_n522_), .O(new_n523_));
  nor2 g0393(.a(new_n235_), .b(i_26_), .O(new_n524_));
  inv1 g0394(.a(new_n524_), .O(new_n525_));
  nor2 g0395(.a(new_n525_), .b(new_n269_), .O(new_n526_));
  inv1 g0396(.a(new_n526_), .O(new_n527_));
  inv1 g0397(.a(i_6_), .O(new_n528_));
  nor2 g0398(.a(new_n528_), .b(i_7_), .O(new_n529_));
  inv1 g0399(.a(new_n529_), .O(new_n530_));
  nor2 g0400(.a(new_n530_), .b(new_n433_), .O(new_n531_));
  inv1 g0401(.a(new_n531_), .O(new_n532_));
  nor2 g0402(.a(new_n161_), .b(i_24_), .O(new_n533_));
  inv1 g0403(.a(new_n533_), .O(new_n534_));
  nor2 g0404(.a(i_11_), .b(i_3_), .O(new_n535_));
  inv1 g0405(.a(new_n535_), .O(new_n536_));
  nor2 g0406(.a(new_n536_), .b(new_n200_), .O(new_n537_));
  inv1 g0407(.a(new_n537_), .O(new_n538_));
  nor2 g0408(.a(new_n538_), .b(new_n534_), .O(new_n539_));
  inv1 g0409(.a(new_n539_), .O(new_n540_));
  nor2 g0410(.a(new_n540_), .b(new_n532_), .O(new_n541_));
  inv1 g0411(.a(new_n541_), .O(new_n542_));
  nor2 g0412(.a(new_n542_), .b(new_n527_), .O(new_n543_));
  inv1 g0413(.a(new_n543_), .O(new_n544_));
  nor2 g0414(.a(new_n544_), .b(new_n523_), .O(o_12_));
  nor2 g0415(.a(new_n286_), .b(i_52_), .O(new_n546_));
  inv1 g0416(.a(new_n546_), .O(new_n547_));
  nor2 g0417(.a(new_n547_), .b(new_n292_), .O(new_n548_));
  inv1 g0418(.a(new_n548_), .O(new_n549_));
  nor2 g0419(.a(new_n271_), .b(i_45_), .O(new_n550_));
  inv1 g0420(.a(new_n550_), .O(new_n551_));
  nor2 g0421(.a(new_n344_), .b(new_n208_), .O(new_n552_));
  inv1 g0422(.a(new_n552_), .O(new_n553_));
  nor2 g0423(.a(new_n553_), .b(new_n551_), .O(new_n554_));
  inv1 g0424(.a(new_n554_), .O(new_n555_));
  nor2 g0425(.a(new_n555_), .b(new_n549_), .O(new_n556_));
  inv1 g0426(.a(new_n556_), .O(new_n557_));
  nor2 g0427(.a(new_n173_), .b(i_51_), .O(new_n558_));
  inv1 g0428(.a(new_n558_), .O(new_n559_));
  nor2 g0429(.a(new_n559_), .b(new_n284_), .O(new_n560_));
  inv1 g0430(.a(new_n560_), .O(new_n561_));
  nor2 g0431(.a(i_37_), .b(i_35_), .O(new_n562_));
  inv1 g0432(.a(new_n562_), .O(new_n563_));
  nor2 g0433(.a(i_60_), .b(i_36_), .O(new_n564_));
  inv1 g0434(.a(new_n564_), .O(new_n565_));
  nor2 g0435(.a(new_n565_), .b(new_n206_), .O(new_n566_));
  inv1 g0436(.a(new_n566_), .O(new_n567_));
  nor2 g0437(.a(new_n567_), .b(new_n563_), .O(new_n568_));
  inv1 g0438(.a(new_n568_), .O(new_n569_));
  nor2 g0439(.a(new_n569_), .b(new_n561_), .O(new_n570_));
  inv1 g0440(.a(new_n570_), .O(new_n571_));
  nor2 g0441(.a(new_n571_), .b(new_n557_), .O(new_n572_));
  inv1 g0442(.a(new_n572_), .O(new_n573_));
  nor2 g0443(.a(new_n327_), .b(new_n253_), .O(new_n574_));
  inv1 g0444(.a(new_n574_), .O(new_n575_));
  inv1 g0445(.a(i_19_), .O(new_n576_));
  nor2 g0446(.a(new_n576_), .b(i_32_), .O(new_n577_));
  inv1 g0447(.a(new_n577_), .O(new_n578_));
  nor2 g0448(.a(new_n578_), .b(new_n145_), .O(new_n579_));
  inv1 g0449(.a(new_n579_), .O(new_n580_));
  nor2 g0450(.a(new_n580_), .b(new_n321_), .O(new_n581_));
  inv1 g0451(.a(new_n581_), .O(new_n582_));
  nor2 g0452(.a(new_n582_), .b(new_n527_), .O(new_n583_));
  inv1 g0453(.a(new_n583_), .O(new_n584_));
  nor2 g0454(.a(new_n584_), .b(new_n575_), .O(new_n585_));
  inv1 g0455(.a(new_n585_), .O(new_n586_));
  nor2 g0456(.a(new_n586_), .b(new_n313_), .O(new_n587_));
  inv1 g0457(.a(new_n587_), .O(new_n588_));
  nor2 g0458(.a(new_n588_), .b(new_n573_), .O(o_37_));
  nor2 g0459(.a(new_n137_), .b(i_22_), .O(new_n590_));
  inv1 g0460(.a(new_n590_), .O(new_n591_));
  nor2 g0461(.a(new_n591_), .b(new_n134_), .O(new_n592_));
  inv1 g0462(.a(new_n592_), .O(new_n593_));
  nor2 g0463(.a(new_n321_), .b(i_21_), .O(new_n594_));
  inv1 g0464(.a(new_n594_), .O(new_n595_));
  nor2 g0465(.a(new_n595_), .b(new_n593_), .O(new_n596_));
  inv1 g0466(.a(new_n596_), .O(new_n597_));
  nor2 g0467(.a(new_n597_), .b(new_n233_), .O(new_n598_));
  inv1 g0468(.a(new_n598_), .O(new_n599_));
  nor2 g0469(.a(i_36_), .b(i_34_), .O(new_n600_));
  inv1 g0470(.a(new_n600_), .O(new_n601_));
  nor2 g0471(.a(new_n601_), .b(i_33_), .O(new_n602_));
  inv1 g0472(.a(new_n602_), .O(new_n603_));
  nor2 g0473(.a(new_n603_), .b(new_n157_), .O(new_n604_));
  inv1 g0474(.a(new_n604_), .O(new_n605_));
  nor2 g0475(.a(new_n393_), .b(i_45_), .O(new_n606_));
  inv1 g0476(.a(new_n606_), .O(new_n607_));
  nor2 g0477(.a(new_n607_), .b(new_n387_), .O(new_n608_));
  inv1 g0478(.a(new_n608_), .O(new_n609_));
  nor2 g0479(.a(new_n609_), .b(new_n605_), .O(new_n610_));
  inv1 g0480(.a(new_n610_), .O(new_n611_));
  nor2 g0481(.a(new_n344_), .b(i_59_), .O(new_n612_));
  inv1 g0482(.a(new_n612_), .O(new_n613_));
  nor2 g0483(.a(new_n613_), .b(new_n210_), .O(new_n614_));
  inv1 g0484(.a(new_n614_), .O(new_n615_));
  nor2 g0485(.a(i_47_), .b(i_49_), .O(new_n616_));
  inv1 g0486(.a(new_n616_), .O(new_n617_));
  nor2 g0487(.a(new_n617_), .b(i_48_), .O(new_n618_));
  inv1 g0488(.a(new_n618_), .O(new_n619_));
  nor2 g0489(.a(new_n190_), .b(i_52_), .O(new_n620_));
  inv1 g0490(.a(new_n620_), .O(new_n621_));
  nor2 g0491(.a(new_n621_), .b(new_n619_), .O(new_n622_));
  inv1 g0492(.a(new_n622_), .O(new_n623_));
  nor2 g0493(.a(new_n623_), .b(new_n615_), .O(new_n624_));
  inv1 g0494(.a(new_n624_), .O(new_n625_));
  nor2 g0495(.a(new_n625_), .b(new_n611_), .O(new_n626_));
  inv1 g0496(.a(new_n626_), .O(new_n627_));
  nor2 g0497(.a(new_n377_), .b(i_57_), .O(new_n628_));
  inv1 g0498(.a(new_n628_), .O(new_n629_));
  nor2 g0499(.a(new_n629_), .b(new_n171_), .O(new_n630_));
  inv1 g0500(.a(new_n630_), .O(new_n631_));
  inv1 g0501(.a(i_32_), .O(new_n632_));
  nor2 g0502(.a(new_n251_), .b(new_n632_), .O(new_n633_));
  inv1 g0503(.a(new_n633_), .O(new_n634_));
  nor2 g0504(.a(new_n634_), .b(new_n631_), .O(new_n635_));
  inv1 g0505(.a(new_n635_), .O(new_n636_));
  nor2 g0506(.a(new_n636_), .b(new_n311_), .O(new_n637_));
  inv1 g0507(.a(new_n637_), .O(new_n638_));
  nor2 g0508(.a(new_n638_), .b(new_n627_), .O(new_n639_));
  inv1 g0509(.a(new_n639_), .O(new_n640_));
  nor2 g0510(.a(new_n640_), .b(new_n599_), .O(o_26_));
  inv1 g0511(.a(i_37_), .O(new_n642_));
  nor2 g0512(.a(new_n501_), .b(new_n642_), .O(o_11_));
  inv1 g0513(.a(i_57_), .O(new_n644_));
  nor2 g0514(.a(new_n186_), .b(new_n644_), .O(new_n645_));
  inv1 g0515(.a(new_n645_), .O(new_n646_));
  nor2 g0516(.a(new_n646_), .b(new_n290_), .O(new_n647_));
  inv1 g0517(.a(new_n647_), .O(new_n648_));
  nor2 g0518(.a(new_n648_), .b(new_n279_), .O(new_n649_));
  inv1 g0519(.a(new_n649_), .O(new_n650_));
  nor2 g0520(.a(new_n650_), .b(new_n263_), .O(o_50_));
  nor2 g0521(.a(new_n200_), .b(i_7_), .O(new_n652_));
  inv1 g0522(.a(new_n652_), .O(new_n653_));
  nor2 g0523(.a(new_n653_), .b(new_n163_), .O(new_n654_));
  inv1 g0524(.a(new_n654_), .O(new_n655_));
  nor2 g0525(.a(i_3_), .b(i_6_), .O(new_n656_));
  inv1 g0526(.a(new_n656_), .O(new_n657_));
  nor2 g0527(.a(new_n657_), .b(i_0_), .O(new_n658_));
  inv1 g0528(.a(new_n658_), .O(new_n659_));
  nor2 g0529(.a(new_n659_), .b(new_n655_), .O(new_n660_));
  inv1 g0530(.a(new_n660_), .O(new_n661_));
  nor2 g0531(.a(new_n267_), .b(i_37_), .O(new_n662_));
  inv1 g0532(.a(new_n662_), .O(new_n663_));
  nor2 g0533(.a(new_n393_), .b(i_41_), .O(new_n664_));
  inv1 g0534(.a(new_n664_), .O(new_n665_));
  nor2 g0535(.a(new_n665_), .b(new_n383_), .O(new_n666_));
  inv1 g0536(.a(new_n666_), .O(new_n667_));
  nor2 g0537(.a(new_n667_), .b(new_n663_), .O(new_n668_));
  inv1 g0538(.a(new_n668_), .O(new_n669_));
  nor2 g0539(.a(new_n669_), .b(new_n661_), .O(new_n670_));
  inv1 g0540(.a(new_n670_), .O(new_n671_));
  nor2 g0541(.a(new_n139_), .b(i_35_), .O(new_n672_));
  inv1 g0542(.a(new_n672_), .O(new_n673_));
  nor2 g0543(.a(new_n673_), .b(new_n241_), .O(new_n674_));
  inv1 g0544(.a(new_n674_), .O(new_n675_));
  inv1 g0545(.a(i_61_), .O(new_n676_));
  nor2 g0546(.a(i_62_), .b(new_n676_), .O(new_n677_));
  inv1 g0547(.a(new_n677_), .O(new_n678_));
  nor2 g0548(.a(new_n678_), .b(new_n471_), .O(new_n679_));
  inv1 g0549(.a(new_n679_), .O(new_n680_));
  nor2 g0550(.a(new_n680_), .b(new_n675_), .O(new_n681_));
  inv1 g0551(.a(new_n681_), .O(new_n682_));
  nor2 g0552(.a(new_n682_), .b(new_n671_), .O(o_36_));
  nor2 g0553(.a(new_n354_), .b(new_n305_), .O(new_n684_));
  inv1 g0554(.a(new_n684_), .O(new_n685_));
  nor2 g0555(.a(new_n685_), .b(new_n368_), .O(new_n686_));
  inv1 g0556(.a(new_n686_), .O(new_n687_));
  nor2 g0557(.a(new_n601_), .b(i_35_), .O(new_n688_));
  inv1 g0558(.a(new_n688_), .O(new_n689_));
  nor2 g0559(.a(new_n689_), .b(new_n275_), .O(new_n690_));
  inv1 g0560(.a(new_n690_), .O(new_n691_));
  inv1 g0561(.a(i_13_), .O(new_n692_));
  nor2 g0562(.a(i_60_), .b(new_n692_), .O(new_n693_));
  inv1 g0563(.a(new_n693_), .O(new_n694_));
  nor2 g0564(.a(new_n694_), .b(new_n307_), .O(new_n695_));
  inv1 g0565(.a(new_n695_), .O(new_n696_));
  nor2 g0566(.a(new_n696_), .b(new_n360_), .O(new_n697_));
  inv1 g0567(.a(new_n697_), .O(new_n698_));
  nor2 g0568(.a(new_n251_), .b(i_33_), .O(new_n699_));
  inv1 g0569(.a(new_n699_), .O(new_n700_));
  nor2 g0570(.a(new_n700_), .b(new_n553_), .O(new_n701_));
  inv1 g0571(.a(new_n701_), .O(new_n702_));
  nor2 g0572(.a(new_n702_), .b(new_n698_), .O(new_n703_));
  inv1 g0573(.a(new_n703_), .O(new_n704_));
  nor2 g0574(.a(new_n704_), .b(new_n691_), .O(new_n705_));
  inv1 g0575(.a(new_n705_), .O(new_n706_));
  nor2 g0576(.a(new_n706_), .b(new_n687_), .O(new_n707_));
  inv1 g0577(.a(new_n707_), .O(new_n708_));
  nor2 g0578(.a(new_n708_), .b(new_n599_), .O(o_27_));
  nor2 g0579(.a(new_n411_), .b(new_n409_), .O(new_n710_));
  inv1 g0580(.a(new_n710_), .O(new_n711_));
  nor2 g0581(.a(new_n711_), .b(i_43_), .O(new_n712_));
  inv1 g0582(.a(new_n712_), .O(new_n713_));
  inv1 g0583(.a(i_50_), .O(new_n714_));
  nor2 g0584(.a(i_58_), .b(new_n714_), .O(new_n715_));
  inv1 g0585(.a(new_n715_), .O(new_n716_));
  nor2 g0586(.a(new_n716_), .b(new_n713_), .O(o_14_));
  nor2 g0587(.a(new_n457_), .b(new_n455_), .O(new_n718_));
  inv1 g0588(.a(new_n718_), .O(new_n719_));
  nor2 g0589(.a(new_n186_), .b(i_51_), .O(new_n720_));
  inv1 g0590(.a(new_n720_), .O(new_n721_));
  nor2 g0591(.a(new_n169_), .b(i_43_), .O(new_n722_));
  inv1 g0592(.a(new_n722_), .O(new_n723_));
  nor2 g0593(.a(new_n723_), .b(new_n721_), .O(new_n724_));
  inv1 g0594(.a(new_n724_), .O(new_n725_));
  nor2 g0595(.a(new_n725_), .b(new_n719_), .O(new_n726_));
  inv1 g0596(.a(new_n726_), .O(new_n727_));
  inv1 g0597(.a(i_4_), .O(new_n728_));
  nor2 g0598(.a(new_n728_), .b(i_3_), .O(new_n729_));
  inv1 g0599(.a(new_n729_), .O(new_n730_));
  nor2 g0600(.a(i_58_), .b(i_0_), .O(new_n731_));
  inv1 g0601(.a(new_n731_), .O(new_n732_));
  nor2 g0602(.a(new_n732_), .b(new_n730_), .O(new_n733_));
  inv1 g0603(.a(new_n733_), .O(new_n734_));
  nor2 g0604(.a(new_n734_), .b(new_n157_), .O(new_n735_));
  inv1 g0605(.a(new_n735_), .O(new_n736_));
  nor2 g0606(.a(new_n437_), .b(new_n210_), .O(new_n737_));
  inv1 g0607(.a(new_n737_), .O(new_n738_));
  nor2 g0608(.a(new_n738_), .b(new_n736_), .O(new_n739_));
  inv1 g0609(.a(new_n739_), .O(new_n740_));
  nor2 g0610(.a(new_n740_), .b(new_n727_), .O(new_n741_));
  inv1 g0611(.a(new_n741_), .O(new_n742_));
  nor2 g0612(.a(new_n742_), .b(new_n465_), .O(o_35_));
  inv1 g0613(.a(i_25_), .O(new_n744_));
  nor2 g0614(.a(new_n435_), .b(i_43_), .O(new_n745_));
  inv1 g0615(.a(new_n745_), .O(new_n746_));
  nor2 g0616(.a(new_n746_), .b(new_n445_), .O(new_n747_));
  inv1 g0617(.a(new_n747_), .O(new_n748_));
  nor2 g0618(.a(new_n748_), .b(new_n744_), .O(new_n749_));
  inv1 g0619(.a(new_n749_), .O(new_n750_));
  nor2 g0620(.a(new_n750_), .b(new_n417_), .O(o_28_));
  nor2 g0621(.a(new_n132_), .b(i_15_), .O(new_n752_));
  inv1 g0622(.a(new_n752_), .O(new_n753_));
  nor2 g0623(.a(new_n753_), .b(new_n455_), .O(new_n754_));
  inv1 g0624(.a(new_n754_), .O(new_n755_));
  nor2 g0625(.a(new_n221_), .b(i_3_), .O(new_n756_));
  inv1 g0626(.a(new_n756_), .O(new_n757_));
  nor2 g0627(.a(new_n757_), .b(new_n755_), .O(new_n758_));
  inv1 g0628(.a(new_n758_), .O(new_n759_));
  nor2 g0629(.a(new_n447_), .b(i_62_), .O(new_n760_));
  inv1 g0630(.a(new_n760_), .O(new_n761_));
  nor2 g0631(.a(new_n155_), .b(i_30_), .O(new_n762_));
  inv1 g0632(.a(new_n762_), .O(new_n763_));
  nor2 g0633(.a(new_n763_), .b(new_n427_), .O(new_n764_));
  inv1 g0634(.a(new_n764_), .O(new_n765_));
  inv1 g0635(.a(i_41_), .O(new_n766_));
  nor2 g0636(.a(new_n766_), .b(i_26_), .O(new_n767_));
  inv1 g0637(.a(new_n767_), .O(new_n768_));
  nor2 g0638(.a(new_n768_), .b(new_n137_), .O(new_n769_));
  inv1 g0639(.a(new_n769_), .O(new_n770_));
  nor2 g0640(.a(new_n770_), .b(new_n437_), .O(new_n771_));
  inv1 g0641(.a(new_n771_), .O(new_n772_));
  nor2 g0642(.a(new_n772_), .b(new_n765_), .O(new_n773_));
  inv1 g0643(.a(new_n773_), .O(new_n774_));
  nor2 g0644(.a(new_n774_), .b(new_n761_), .O(new_n775_));
  inv1 g0645(.a(new_n775_), .O(new_n776_));
  nor2 g0646(.a(new_n776_), .b(new_n759_), .O(o_13_));
  inv1 g0647(.a(i_58_), .O(new_n778_));
  nor2 g0648(.a(new_n413_), .b(new_n161_), .O(new_n779_));
  inv1 g0649(.a(new_n779_), .O(new_n780_));
  nor2 g0650(.a(new_n780_), .b(new_n778_), .O(o_34_));
  nor2 g0651(.a(new_n433_), .b(new_n241_), .O(new_n782_));
  inv1 g0652(.a(new_n782_), .O(new_n783_));
  nor2 g0653(.a(new_n783_), .b(new_n521_), .O(new_n784_));
  inv1 g0654(.a(new_n784_), .O(new_n785_));
  nor2 g0655(.a(new_n269_), .b(new_n175_), .O(new_n786_));
  inv1 g0656(.a(new_n786_), .O(new_n787_));
  inv1 g0657(.a(i_0_), .O(new_n788_));
  nor2 g0658(.a(new_n657_), .b(new_n788_), .O(new_n789_));
  inv1 g0659(.a(new_n789_), .O(new_n790_));
  nor2 g0660(.a(new_n790_), .b(new_n655_), .O(new_n791_));
  inv1 g0661(.a(new_n791_), .O(new_n792_));
  nor2 g0662(.a(new_n792_), .b(new_n787_), .O(new_n793_));
  inv1 g0663(.a(new_n793_), .O(new_n794_));
  nor2 g0664(.a(new_n794_), .b(new_n785_), .O(o_21_));
  nor2 g0665(.a(new_n521_), .b(i_47_), .O(new_n796_));
  inv1 g0666(.a(new_n796_), .O(new_n797_));
  nor2 g0667(.a(new_n765_), .b(i_46_), .O(new_n798_));
  inv1 g0668(.a(new_n798_), .O(new_n799_));
  inv1 g0669(.a(i_26_), .O(new_n800_));
  nor2 g0670(.a(new_n137_), .b(new_n800_), .O(new_n801_));
  inv1 g0671(.a(new_n801_), .O(new_n802_));
  nor2 g0672(.a(new_n802_), .b(new_n759_), .O(new_n803_));
  inv1 g0673(.a(new_n803_), .O(new_n804_));
  nor2 g0674(.a(new_n804_), .b(new_n799_), .O(new_n805_));
  inv1 g0675(.a(new_n805_), .O(new_n806_));
  nor2 g0676(.a(new_n806_), .b(new_n797_), .O(o_16_));
  nor2 g0677(.a(new_n459_), .b(new_n249_), .O(new_n808_));
  inv1 g0678(.a(new_n808_), .O(new_n809_));
  nor2 g0679(.a(new_n809_), .b(new_n245_), .O(new_n810_));
  inv1 g0680(.a(new_n810_), .O(new_n811_));
  nor2 g0681(.a(new_n563_), .b(i_34_), .O(new_n812_));
  inv1 g0682(.a(new_n812_), .O(new_n813_));
  nor2 g0683(.a(new_n813_), .b(new_n269_), .O(new_n814_));
  inv1 g0684(.a(new_n814_), .O(new_n815_));
  nor2 g0685(.a(new_n139_), .b(i_33_), .O(new_n816_));
  inv1 g0686(.a(new_n816_), .O(new_n817_));
  nor2 g0687(.a(new_n817_), .b(new_n815_), .O(new_n818_));
  inv1 g0688(.a(new_n818_), .O(new_n819_));
  nor2 g0689(.a(new_n819_), .b(new_n811_), .O(new_n820_));
  inv1 g0690(.a(new_n820_), .O(new_n821_));
  nor2 g0691(.a(new_n393_), .b(i_42_), .O(new_n822_));
  inv1 g0692(.a(new_n822_), .O(new_n823_));
  nor2 g0693(.a(new_n823_), .b(new_n383_), .O(new_n824_));
  inv1 g0694(.a(new_n824_), .O(new_n825_));
  nor2 g0695(.a(new_n825_), .b(new_n212_), .O(new_n826_));
  inv1 g0696(.a(new_n826_), .O(new_n827_));
  inv1 g0697(.a(i_54_), .O(new_n828_));
  nor2 g0698(.a(new_n186_), .b(new_n828_), .O(new_n829_));
  inv1 g0699(.a(new_n829_), .O(new_n830_));
  nor2 g0700(.a(new_n830_), .b(new_n827_), .O(new_n831_));
  inv1 g0701(.a(new_n831_), .O(new_n832_));
  nor2 g0702(.a(new_n832_), .b(new_n821_), .O(o_40_));
  inv1 g0703(.a(i_39_), .O(new_n834_));
  nor2 g0704(.a(new_n420_), .b(new_n834_), .O(new_n835_));
  inv1 g0705(.a(new_n835_), .O(new_n836_));
  nor2 g0706(.a(new_n836_), .b(new_n427_), .O(new_n837_));
  inv1 g0707(.a(new_n837_), .O(new_n838_));
  nor2 g0708(.a(new_n838_), .b(new_n711_), .O(o_33_));
  nor2 g0709(.a(new_n233_), .b(new_n149_), .O(new_n840_));
  inv1 g0710(.a(new_n840_), .O(new_n841_));
  inv1 g0711(.a(i_36_), .O(new_n842_));
  nor2 g0712(.a(new_n563_), .b(new_n842_), .O(new_n843_));
  inv1 g0713(.a(new_n843_), .O(new_n844_));
  nor2 g0714(.a(new_n844_), .b(new_n153_), .O(new_n845_));
  inv1 g0715(.a(new_n845_), .O(new_n846_));
  nor2 g0716(.a(new_n269_), .b(new_n249_), .O(new_n847_));
  inv1 g0717(.a(new_n847_), .O(new_n848_));
  nor2 g0718(.a(new_n848_), .b(new_n846_), .O(new_n849_));
  inv1 g0719(.a(new_n849_), .O(new_n850_));
  nor2 g0720(.a(new_n850_), .b(new_n561_), .O(new_n851_));
  inv1 g0721(.a(new_n851_), .O(new_n852_));
  nor2 g0722(.a(new_n629_), .b(new_n615_), .O(new_n853_));
  inv1 g0723(.a(new_n853_), .O(new_n854_));
  nor2 g0724(.a(new_n161_), .b(i_12_), .O(new_n855_));
  inv1 g0725(.a(new_n855_), .O(new_n856_));
  nor2 g0726(.a(new_n551_), .b(new_n387_), .O(new_n857_));
  inv1 g0727(.a(new_n857_), .O(new_n858_));
  nor2 g0728(.a(new_n858_), .b(new_n856_), .O(new_n859_));
  inv1 g0729(.a(new_n859_), .O(new_n860_));
  nor2 g0730(.a(new_n860_), .b(new_n854_), .O(new_n861_));
  inv1 g0731(.a(new_n861_), .O(new_n862_));
  nor2 g0732(.a(new_n862_), .b(new_n852_), .O(new_n863_));
  inv1 g0733(.a(new_n863_), .O(new_n864_));
  nor2 g0734(.a(new_n864_), .b(new_n841_), .O(o_22_));
  inv1 g0735(.a(i_10_), .O(new_n866_));
  nor2 g0736(.a(i_58_), .b(new_n866_), .O(new_n867_));
  inv1 g0737(.a(new_n867_), .O(new_n868_));
  nor2 g0738(.a(new_n868_), .b(new_n780_), .O(o_15_));
  inv1 g0739(.a(i_46_), .O(new_n870_));
  nor2 g0740(.a(new_n420_), .b(new_n870_), .O(new_n871_));
  inv1 g0741(.a(new_n871_), .O(new_n872_));
  nor2 g0742(.a(new_n872_), .b(new_n417_), .O(o_32_));
  inv1 g0743(.a(i_16_), .O(new_n874_));
  nor2 g0744(.a(i_17_), .b(i_18_), .O(new_n875_));
  inv1 g0745(.a(new_n875_), .O(new_n876_));
  nor2 g0746(.a(new_n876_), .b(new_n874_), .O(new_n877_));
  inv1 g0747(.a(new_n877_), .O(new_n878_));
  nor2 g0748(.a(new_n878_), .b(new_n525_), .O(new_n879_));
  inv1 g0749(.a(new_n879_), .O(new_n880_));
  nor2 g0750(.a(new_n880_), .b(new_n575_), .O(new_n881_));
  inv1 g0751(.a(new_n881_), .O(new_n882_));
  nor2 g0752(.a(new_n856_), .b(new_n249_), .O(new_n883_));
  inv1 g0753(.a(new_n883_), .O(new_n884_));
  nor2 g0754(.a(new_n884_), .b(new_n631_), .O(new_n885_));
  inv1 g0755(.a(new_n885_), .O(new_n886_));
  nor2 g0756(.a(new_n886_), .b(new_n882_), .O(new_n887_));
  inv1 g0757(.a(new_n887_), .O(new_n888_));
  nor2 g0758(.a(new_n888_), .b(new_n233_), .O(new_n889_));
  inv1 g0759(.a(new_n889_), .O(new_n890_));
  nor2 g0760(.a(new_n890_), .b(new_n627_), .O(o_23_));
  inv1 g0761(.a(i_62_), .O(new_n892_));
  nor2 g0762(.a(new_n447_), .b(new_n892_), .O(new_n893_));
  inv1 g0763(.a(new_n893_), .O(new_n894_));
  nor2 g0764(.a(new_n894_), .b(new_n653_), .O(new_n895_));
  inv1 g0765(.a(new_n895_), .O(new_n896_));
  nor2 g0766(.a(new_n896_), .b(new_n443_), .O(o_18_));
  nor2 g0767(.a(new_n700_), .b(new_n593_), .O(new_n898_));
  inv1 g0768(.a(new_n898_), .O(new_n899_));
  nor2 g0769(.a(new_n899_), .b(new_n233_), .O(new_n900_));
  inv1 g0770(.a(new_n900_), .O(new_n901_));
  nor2 g0771(.a(new_n876_), .b(i_64_), .O(new_n902_));
  inv1 g0772(.a(new_n902_), .O(new_n903_));
  inv1 g0773(.a(i_21_), .O(new_n904_));
  nor2 g0774(.a(new_n265_), .b(new_n904_), .O(new_n905_));
  inv1 g0775(.a(new_n905_), .O(new_n906_));
  nor2 g0776(.a(new_n906_), .b(new_n903_), .O(new_n907_));
  inv1 g0777(.a(new_n907_), .O(new_n908_));
  nor2 g0778(.a(new_n884_), .b(new_n290_), .O(new_n909_));
  inv1 g0779(.a(new_n909_), .O(new_n910_));
  nor2 g0780(.a(new_n910_), .b(new_n908_), .O(new_n911_));
  inv1 g0781(.a(new_n911_), .O(new_n912_));
  nor2 g0782(.a(new_n292_), .b(i_63_), .O(new_n913_));
  inv1 g0783(.a(new_n913_), .O(new_n914_));
  nor2 g0784(.a(new_n914_), .b(new_n212_), .O(new_n915_));
  inv1 g0785(.a(new_n915_), .O(new_n916_));
  nor2 g0786(.a(new_n916_), .b(new_n691_), .O(new_n917_));
  inv1 g0787(.a(new_n917_), .O(new_n918_));
  nor2 g0788(.a(new_n918_), .b(new_n912_), .O(new_n919_));
  inv1 g0789(.a(new_n919_), .O(new_n920_));
  nor2 g0790(.a(new_n920_), .b(new_n901_), .O(o_31_));
  inv1 g0791(.a(i_11_), .O(new_n922_));
  nor2 g0792(.a(i_60_), .b(new_n922_), .O(new_n923_));
  inv1 g0793(.a(new_n923_), .O(new_n924_));
  nor2 g0794(.a(new_n924_), .b(new_n503_), .O(new_n925_));
  inv1 g0795(.a(new_n925_), .O(new_n926_));
  nor2 g0796(.a(new_n926_), .b(new_n422_), .O(new_n927_));
  inv1 g0797(.a(new_n927_), .O(new_n928_));
  nor2 g0798(.a(new_n928_), .b(new_n753_), .O(new_n929_));
  inv1 g0799(.a(new_n929_), .O(new_n930_));
  nor2 g0800(.a(new_n930_), .b(new_n415_), .O(o_24_));
  nor2 g0801(.a(new_n663_), .b(new_n141_), .O(new_n932_));
  inv1 g0802(.a(new_n932_), .O(new_n933_));
  nor2 g0803(.a(new_n933_), .b(new_n755_), .O(new_n934_));
  inv1 g0804(.a(new_n934_), .O(new_n935_));
  inv1 g0805(.a(i_3_), .O(new_n936_));
  nor2 g0806(.a(new_n221_), .b(new_n936_), .O(new_n937_));
  inv1 g0807(.a(new_n937_), .O(new_n938_));
  nor2 g0808(.a(new_n938_), .b(new_n935_), .O(new_n939_));
  inv1 g0809(.a(new_n939_), .O(new_n940_));
  nor2 g0810(.a(new_n940_), .b(new_n523_), .O(o_17_));
  inv1 g0811(.a(i_20_), .O(new_n942_));
  nor2 g0812(.a(i_21_), .b(new_n942_), .O(new_n943_));
  inv1 g0813(.a(new_n943_), .O(new_n944_));
  nor2 g0814(.a(new_n944_), .b(i_16_), .O(new_n945_));
  inv1 g0815(.a(new_n945_), .O(new_n946_));
  nor2 g0816(.a(new_n946_), .b(new_n153_), .O(new_n947_));
  inv1 g0817(.a(new_n947_), .O(new_n948_));
  nor2 g0818(.a(new_n948_), .b(new_n269_), .O(new_n949_));
  inv1 g0819(.a(new_n949_), .O(new_n950_));
  nor2 g0820(.a(new_n950_), .b(new_n884_), .O(new_n951_));
  inv1 g0821(.a(new_n951_), .O(new_n952_));
  nor2 g0822(.a(new_n952_), .b(new_n573_), .O(new_n953_));
  inv1 g0823(.a(new_n953_), .O(new_n954_));
  nor2 g0824(.a(new_n954_), .b(new_n841_), .O(o_56_));
  inv1 g0825(.a(i_1_), .O(new_n956_));
  nor2 g0826(.a(i_2_), .b(new_n956_), .O(new_n957_));
  inv1 g0827(.a(new_n957_), .O(new_n958_));
  nor2 g0828(.a(new_n958_), .b(i_0_), .O(new_n959_));
  inv1 g0829(.a(new_n959_), .O(new_n960_));
  nor2 g0830(.a(new_n960_), .b(new_n194_), .O(new_n961_));
  inv1 g0831(.a(new_n961_), .O(new_n962_));
  nor2 g0832(.a(new_n962_), .b(new_n227_), .O(new_n963_));
  inv1 g0833(.a(new_n963_), .O(new_n964_));
  nor2 g0834(.a(new_n964_), .b(new_n261_), .O(new_n965_));
  inv1 g0835(.a(new_n965_), .O(new_n966_));
  nor2 g0836(.a(new_n966_), .b(new_n279_), .O(o_43_));
  nor2 g0837(.a(new_n362_), .b(new_n354_), .O(new_n968_));
  inv1 g0838(.a(new_n968_), .O(new_n969_));
  nor2 g0839(.a(new_n969_), .b(new_n884_), .O(new_n970_));
  inv1 g0840(.a(new_n970_), .O(new_n971_));
  nor2 g0841(.a(i_21_), .b(i_63_), .O(new_n972_));
  inv1 g0842(.a(new_n972_), .O(new_n973_));
  inv1 g0843(.a(i_52_), .O(new_n974_));
  nor2 g0844(.a(new_n974_), .b(i_53_), .O(new_n975_));
  inv1 g0845(.a(new_n975_), .O(new_n976_));
  nor2 g0846(.a(new_n976_), .b(i_51_), .O(new_n977_));
  inv1 g0847(.a(new_n977_), .O(new_n978_));
  nor2 g0848(.a(new_n978_), .b(new_n973_), .O(new_n979_));
  inv1 g0849(.a(new_n979_), .O(new_n980_));
  nor2 g0850(.a(new_n903_), .b(new_n188_), .O(new_n981_));
  inv1 g0851(.a(new_n981_), .O(new_n982_));
  nor2 g0852(.a(new_n982_), .b(new_n980_), .O(new_n983_));
  inv1 g0853(.a(new_n983_), .O(new_n984_));
  nor2 g0854(.a(new_n984_), .b(new_n691_), .O(new_n985_));
  inv1 g0855(.a(new_n985_), .O(new_n986_));
  nor2 g0856(.a(new_n986_), .b(new_n971_), .O(new_n987_));
  inv1 g0857(.a(new_n987_), .O(new_n988_));
  nor2 g0858(.a(new_n988_), .b(new_n901_), .O(o_30_));
  nor2 g0859(.a(new_n761_), .b(new_n671_), .O(new_n990_));
  inv1 g0860(.a(new_n990_), .O(new_n991_));
  inv1 g0861(.a(i_35_), .O(new_n992_));
  nor2 g0862(.a(new_n139_), .b(new_n992_), .O(new_n993_));
  inv1 g0863(.a(new_n993_), .O(new_n994_));
  nor2 g0864(.a(new_n994_), .b(new_n241_), .O(new_n995_));
  inv1 g0865(.a(new_n995_), .O(new_n996_));
  nor2 g0866(.a(new_n996_), .b(new_n991_), .O(o_55_));
  nor2 g0867(.a(i_9_), .b(i_62_), .O(new_n998_));
  inv1 g0868(.a(new_n998_), .O(new_n999_));
  nor2 g0869(.a(new_n999_), .b(new_n221_), .O(new_n1000_));
  inv1 g0870(.a(new_n1000_), .O(new_n1001_));
  nor2 g0871(.a(new_n1001_), .b(new_n876_), .O(new_n1002_));
  inv1 g0872(.a(new_n1002_), .O(new_n1003_));
  inv1 g0873(.a(i_2_), .O(new_n1004_));
  nor2 g0874(.a(i_0_), .b(new_n1004_), .O(new_n1005_));
  inv1 g0875(.a(new_n1005_), .O(new_n1006_));
  nor2 g0876(.a(new_n1006_), .b(i_15_), .O(new_n1007_));
  inv1 g0877(.a(new_n1007_), .O(new_n1008_));
  nor2 g0878(.a(new_n1008_), .b(new_n225_), .O(new_n1009_));
  inv1 g0879(.a(new_n1009_), .O(new_n1010_));
  nor2 g0880(.a(new_n1010_), .b(new_n1003_), .O(new_n1011_));
  inv1 g0881(.a(new_n1011_), .O(new_n1012_));
  nor2 g0882(.a(i_59_), .b(i_61_), .O(new_n1013_));
  inv1 g0883(.a(new_n1013_), .O(new_n1014_));
  nor2 g0884(.a(new_n1014_), .b(new_n471_), .O(new_n1015_));
  inv1 g0885(.a(new_n1015_), .O(new_n1016_));
  nor2 g0886(.a(new_n1016_), .b(new_n815_), .O(new_n1017_));
  inv1 g0887(.a(new_n1017_), .O(new_n1018_));
  nor2 g0888(.a(new_n1018_), .b(new_n1012_), .O(new_n1019_));
  inv1 g0889(.a(new_n1019_), .O(new_n1020_));
  nor2 g0890(.a(new_n437_), .b(new_n288_), .O(new_n1021_));
  inv1 g0891(.a(new_n1021_), .O(new_n1022_));
  nor2 g0892(.a(new_n551_), .b(new_n455_), .O(new_n1023_));
  inv1 g0893(.a(new_n1023_), .O(new_n1024_));
  nor2 g0894(.a(new_n1024_), .b(new_n1022_), .O(new_n1025_));
  inv1 g0895(.a(new_n1025_), .O(new_n1026_));
  nor2 g0896(.a(new_n1026_), .b(new_n899_), .O(new_n1027_));
  inv1 g0897(.a(new_n1027_), .O(new_n1028_));
  nor2 g0898(.a(new_n1028_), .b(new_n1020_), .O(o_44_));
  inv1 g0899(.a(i_22_), .O(new_n1030_));
  nor2 g0900(.a(new_n161_), .b(new_n1030_), .O(new_n1031_));
  inv1 g0901(.a(new_n1031_), .O(new_n1032_));
  nor2 g0902(.a(new_n1032_), .b(new_n665_), .O(new_n1033_));
  inv1 g0903(.a(new_n1033_), .O(new_n1034_));
  nor2 g0904(.a(new_n1034_), .b(new_n663_), .O(new_n1035_));
  inv1 g0905(.a(new_n1035_), .O(new_n1036_));
  nor2 g0906(.a(new_n538_), .b(new_n178_), .O(new_n1037_));
  inv1 g0907(.a(new_n1037_), .O(new_n1038_));
  nor2 g0908(.a(new_n1038_), .b(new_n143_), .O(new_n1039_));
  inv1 g0909(.a(new_n1039_), .O(new_n1040_));
  nor2 g0910(.a(new_n1040_), .b(new_n1036_), .O(new_n1041_));
  inv1 g0911(.a(new_n1041_), .O(new_n1042_));
  nor2 g0912(.a(new_n1042_), .b(new_n797_), .O(o_58_));
  inv1 g0913(.a(i_33_), .O(new_n1044_));
  nor2 g0914(.a(new_n139_), .b(new_n1044_), .O(new_n1045_));
  inv1 g0915(.a(new_n1045_), .O(new_n1046_));
  nor2 g0916(.a(new_n1046_), .b(new_n383_), .O(new_n1047_));
  inv1 g0917(.a(new_n1047_), .O(new_n1048_));
  nor2 g0918(.a(new_n377_), .b(i_55_), .O(new_n1049_));
  inv1 g0919(.a(new_n1049_), .O(new_n1050_));
  nor2 g0920(.a(new_n1050_), .b(new_n823_), .O(new_n1051_));
  inv1 g0921(.a(new_n1051_), .O(new_n1052_));
  nor2 g0922(.a(new_n1052_), .b(new_n1048_), .O(new_n1053_));
  inv1 g0923(.a(new_n1053_), .O(new_n1054_));
  nor2 g0924(.a(new_n815_), .b(new_n379_), .O(new_n1055_));
  inv1 g0925(.a(new_n1055_), .O(new_n1056_));
  nor2 g0926(.a(new_n1056_), .b(new_n1054_), .O(new_n1057_));
  inv1 g0927(.a(new_n1057_), .O(new_n1058_));
  nor2 g0928(.a(new_n1058_), .b(new_n811_), .O(o_41_));
  inv1 g0929(.a(i_18_), .O(new_n1060_));
  nor2 g0930(.a(new_n161_), .b(new_n1060_), .O(new_n1061_));
  inv1 g0931(.a(new_n1061_), .O(new_n1062_));
  nor2 g0932(.a(new_n1062_), .b(new_n437_), .O(new_n1063_));
  inv1 g0933(.a(new_n1063_), .O(new_n1064_));
  nor2 g0934(.a(new_n763_), .b(new_n723_), .O(new_n1065_));
  inv1 g0935(.a(new_n1065_), .O(new_n1066_));
  nor2 g0936(.a(new_n1066_), .b(new_n1064_), .O(new_n1067_));
  inv1 g0937(.a(new_n1067_), .O(new_n1068_));
  nor2 g0938(.a(new_n761_), .b(new_n593_), .O(new_n1069_));
  inv1 g0939(.a(new_n1069_), .O(new_n1070_));
  nor2 g0940(.a(new_n1070_), .b(new_n1038_), .O(new_n1071_));
  inv1 g0941(.a(new_n1071_), .O(new_n1072_));
  nor2 g0942(.a(new_n1072_), .b(new_n1068_), .O(o_57_));
  inv1 g0943(.a(i_49_), .O(new_n1074_));
  nor2 g0944(.a(new_n190_), .b(new_n1074_), .O(new_n1075_));
  inv1 g0945(.a(new_n1075_), .O(new_n1076_));
  nor2 g0946(.a(new_n1076_), .b(new_n387_), .O(new_n1077_));
  inv1 g0947(.a(new_n1077_), .O(new_n1078_));
  nor2 g0948(.a(new_n1078_), .b(new_n277_), .O(new_n1079_));
  inv1 g0949(.a(new_n1079_), .O(new_n1080_));
  nor2 g0950(.a(new_n1080_), .b(new_n381_), .O(new_n1081_));
  inv1 g0951(.a(new_n1081_), .O(new_n1082_));
  nor2 g0952(.a(new_n1082_), .b(new_n263_), .O(o_42_));
  inv1 g0953(.a(i_51_), .O(new_n1084_));
  nor2 g0954(.a(new_n787_), .b(new_n1084_), .O(new_n1085_));
  inv1 g0955(.a(new_n1085_), .O(new_n1086_));
  nor2 g0956(.a(new_n1086_), .b(new_n661_), .O(new_n1087_));
  inv1 g0957(.a(new_n1087_), .O(new_n1088_));
  nor2 g0958(.a(new_n1088_), .b(new_n785_), .O(o_20_));
  nor2 g0959(.a(new_n607_), .b(new_n171_), .O(new_n1090_));
  inv1 g0960(.a(new_n1090_), .O(new_n1091_));
  inv1 g0961(.a(i_12_), .O(new_n1092_));
  nor2 g0962(.a(new_n161_), .b(new_n1092_), .O(new_n1093_));
  inv1 g0963(.a(new_n1093_), .O(new_n1094_));
  nor2 g0964(.a(new_n1094_), .b(new_n188_), .O(new_n1095_));
  inv1 g0965(.a(new_n1095_), .O(new_n1096_));
  nor2 g0966(.a(new_n1096_), .b(new_n159_), .O(new_n1097_));
  inv1 g0967(.a(new_n1097_), .O(new_n1098_));
  nor2 g0968(.a(new_n1098_), .b(new_n1091_), .O(new_n1099_));
  inv1 g0969(.a(new_n1099_), .O(new_n1100_));
  nor2 g0970(.a(new_n362_), .b(new_n344_), .O(new_n1101_));
  inv1 g0971(.a(new_n1101_), .O(new_n1102_));
  nor2 g0972(.a(new_n249_), .b(new_n192_), .O(new_n1103_));
  inv1 g0973(.a(new_n1103_), .O(new_n1104_));
  nor2 g0974(.a(new_n1104_), .b(new_n619_), .O(new_n1105_));
  inv1 g0975(.a(new_n1105_), .O(new_n1106_));
  nor2 g0976(.a(new_n1106_), .b(new_n1102_), .O(new_n1107_));
  inv1 g0977(.a(new_n1107_), .O(new_n1108_));
  nor2 g0978(.a(new_n1108_), .b(new_n1100_), .O(new_n1109_));
  inv1 g0979(.a(new_n1109_), .O(new_n1110_));
  nor2 g0980(.a(new_n1110_), .b(new_n841_), .O(o_52_));
  nor2 g0981(.a(new_n825_), .b(new_n241_), .O(new_n1112_));
  inv1 g0982(.a(new_n1112_), .O(new_n1113_));
  nor2 g0983(.a(new_n1113_), .b(new_n1016_), .O(new_n1114_));
  inv1 g0984(.a(new_n1114_), .O(new_n1115_));
  inv1 g0985(.a(i_17_), .O(new_n1116_));
  nor2 g0986(.a(i_30_), .b(i_62_), .O(new_n1117_));
  inv1 g0987(.a(new_n1117_), .O(new_n1118_));
  nor2 g0988(.a(new_n1118_), .b(new_n1116_), .O(new_n1119_));
  inv1 g0989(.a(new_n1119_), .O(new_n1120_));
  nor2 g0990(.a(new_n563_), .b(new_n501_), .O(new_n1121_));
  inv1 g0991(.a(new_n1121_), .O(new_n1122_));
  nor2 g0992(.a(new_n1122_), .b(new_n1120_), .O(new_n1123_));
  inv1 g0993(.a(new_n1123_), .O(new_n1124_));
  nor2 g0994(.a(new_n1124_), .b(new_n269_), .O(new_n1125_));
  inv1 g0995(.a(new_n1125_), .O(new_n1126_));
  nor2 g0996(.a(new_n1126_), .b(new_n461_), .O(new_n1127_));
  inv1 g0997(.a(new_n1127_), .O(new_n1128_));
  nor2 g0998(.a(new_n1128_), .b(new_n1115_), .O(o_47_));
  nor2 g0999(.a(new_n379_), .b(new_n275_), .O(new_n1130_));
  inv1 g1000(.a(new_n1130_), .O(new_n1131_));
  nor2 g1001(.a(new_n1050_), .b(new_n288_), .O(new_n1132_));
  inv1 g1002(.a(new_n1132_), .O(new_n1133_));
  inv1 g1003(.a(i_48_), .O(new_n1134_));
  nor2 g1004(.a(new_n282_), .b(new_n1134_), .O(new_n1135_));
  inv1 g1005(.a(new_n1135_), .O(new_n1136_));
  nor2 g1006(.a(new_n1136_), .b(new_n265_), .O(new_n1137_));
  inv1 g1007(.a(new_n1137_), .O(new_n1138_));
  nor2 g1008(.a(new_n1138_), .b(new_n1133_), .O(new_n1139_));
  inv1 g1009(.a(new_n1139_), .O(new_n1140_));
  nor2 g1010(.a(new_n1140_), .b(new_n1131_), .O(new_n1141_));
  inv1 g1011(.a(new_n1141_), .O(new_n1142_));
  nor2 g1012(.a(new_n1142_), .b(new_n263_), .O(o_51_));
  nor2 g1013(.a(new_n673_), .b(new_n437_), .O(new_n1144_));
  inv1 g1014(.a(new_n1144_), .O(new_n1145_));
  inv1 g1015(.a(i_31_), .O(new_n1146_));
  nor2 g1016(.a(new_n145_), .b(new_n1146_), .O(new_n1147_));
  inv1 g1017(.a(new_n1147_), .O(new_n1148_));
  nor2 g1018(.a(new_n1148_), .b(new_n1133_), .O(new_n1149_));
  inv1 g1019(.a(new_n1149_), .O(new_n1150_));
  nor2 g1020(.a(new_n1150_), .b(new_n1145_), .O(new_n1151_));
  inv1 g1021(.a(new_n1151_), .O(new_n1152_));
  nor2 g1022(.a(new_n1152_), .b(new_n1131_), .O(new_n1153_));
  inv1 g1023(.a(new_n1153_), .O(new_n1154_));
  nor2 g1024(.a(new_n1154_), .b(new_n811_), .O(o_48_));
  inv1 g1025(.a(i_55_), .O(new_n1156_));
  nor2 g1026(.a(new_n675_), .b(new_n1156_), .O(new_n1157_));
  inv1 g1027(.a(new_n1157_), .O(new_n1158_));
  nor2 g1028(.a(new_n1158_), .b(new_n991_), .O(o_54_));
  inv1 g1029(.a(i_34_), .O(new_n1160_));
  nor2 g1030(.a(new_n139_), .b(new_n1160_), .O(new_n1161_));
  inv1 g1031(.a(new_n1161_), .O(new_n1162_));
  nor2 g1032(.a(new_n1162_), .b(new_n469_), .O(new_n1163_));
  inv1 g1033(.a(new_n1163_), .O(new_n1164_));
  nor2 g1034(.a(new_n1164_), .b(new_n487_), .O(new_n1165_));
  inv1 g1035(.a(new_n1165_), .O(new_n1166_));
  nor2 g1036(.a(new_n1166_), .b(new_n381_), .O(new_n1167_));
  inv1 g1037(.a(new_n1167_), .O(new_n1168_));
  nor2 g1038(.a(new_n1168_), .b(new_n811_), .O(o_45_));
  inv1 g1039(.a(i_28_), .O(new_n1170_));
  nor2 g1040(.a(i_37_), .b(new_n1170_), .O(new_n1171_));
  inv1 g1041(.a(new_n1171_), .O(new_n1172_));
  nor2 g1042(.a(new_n1172_), .b(new_n501_), .O(o_10_));
  inv1 g1043(.a(i_63_), .O(new_n1174_));
  nor2 g1044(.a(i_64_), .b(new_n1174_), .O(new_n1175_));
  inv1 g1045(.a(new_n1175_), .O(new_n1176_));
  nor2 g1046(.a(new_n1176_), .b(new_n212_), .O(new_n1177_));
  inv1 g1047(.a(new_n1177_), .O(new_n1178_));
  nor2 g1048(.a(new_n1178_), .b(new_n277_), .O(new_n1179_));
  inv1 g1049(.a(new_n1179_), .O(new_n1180_));
  nor2 g1050(.a(new_n1180_), .b(new_n294_), .O(new_n1181_));
  inv1 g1051(.a(new_n1181_), .O(new_n1182_));
  nor2 g1052(.a(new_n1182_), .b(new_n263_), .O(o_53_));
  nor2 g1053(.a(new_n459_), .b(new_n275_), .O(new_n1184_));
  inv1 g1054(.a(new_n1184_), .O(new_n1185_));
  nor2 g1055(.a(new_n1185_), .b(new_n1145_), .O(new_n1186_));
  inv1 g1056(.a(new_n1186_), .O(new_n1187_));
  inv1 g1057(.a(i_9_), .O(new_n1188_));
  nor2 g1058(.a(new_n247_), .b(new_n1188_), .O(new_n1189_));
  inv1 g1059(.a(new_n1189_), .O(new_n1190_));
  nor2 g1060(.a(new_n1190_), .b(new_n721_), .O(new_n1191_));
  inv1 g1061(.a(new_n1191_), .O(new_n1192_));
  nor2 g1062(.a(new_n1192_), .b(new_n212_), .O(new_n1193_));
  inv1 g1063(.a(new_n1193_), .O(new_n1194_));
  nor2 g1064(.a(new_n1194_), .b(new_n245_), .O(new_n1195_));
  inv1 g1065(.a(new_n1195_), .O(new_n1196_));
  nor2 g1066(.a(new_n1196_), .b(new_n1187_), .O(o_46_));
  inv1 g1067(.a(i_8_), .O(new_n1198_));
  nor2 g1068(.a(i_47_), .b(new_n1198_), .O(new_n1199_));
  inv1 g1069(.a(new_n1199_), .O(new_n1200_));
  nor2 g1070(.a(new_n1200_), .b(new_n135_), .O(new_n1201_));
  inv1 g1071(.a(new_n1201_), .O(new_n1202_));
  nor2 g1072(.a(new_n247_), .b(new_n235_), .O(new_n1203_));
  inv1 g1073(.a(new_n1203_), .O(new_n1204_));
  nor2 g1074(.a(new_n1204_), .b(new_n1202_), .O(new_n1205_));
  inv1 g1075(.a(new_n1205_), .O(new_n1206_));
  nor2 g1076(.a(new_n1206_), .b(new_n534_), .O(new_n1207_));
  inv1 g1077(.a(new_n1207_), .O(new_n1208_));
  nor2 g1078(.a(new_n1208_), .b(new_n519_), .O(new_n1209_));
  inv1 g1079(.a(new_n1209_), .O(new_n1210_));
  nor2 g1080(.a(new_n1210_), .b(new_n799_), .O(o_61_));
  nor2 g1081(.a(new_n346_), .b(i_32_), .O(new_n1212_));
  inv1 g1082(.a(new_n1212_), .O(new_n1213_));
  nor2 g1083(.a(new_n1213_), .b(new_n356_), .O(new_n1214_));
  inv1 g1084(.a(new_n1214_), .O(new_n1215_));
  nor2 g1085(.a(new_n1102_), .b(new_n277_), .O(new_n1216_));
  inv1 g1086(.a(new_n1216_), .O(new_n1217_));
  nor2 g1087(.a(new_n1217_), .b(new_n1215_), .O(new_n1218_));
  inv1 g1088(.a(new_n1218_), .O(new_n1219_));
  inv1 g1089(.a(new_n319_), .O(new_n1220_));
  nor2 g1090(.a(new_n323_), .b(new_n284_), .O(new_n1221_));
  inv1 g1091(.a(new_n1221_), .O(new_n1222_));
  nor2 g1092(.a(new_n1222_), .b(new_n1220_), .O(new_n1223_));
  inv1 g1093(.a(new_n1223_), .O(new_n1224_));
  nor2 g1094(.a(new_n1224_), .b(new_n368_), .O(new_n1225_));
  inv1 g1095(.a(new_n1225_), .O(new_n1226_));
  nor2 g1096(.a(new_n1226_), .b(new_n313_), .O(new_n1227_));
  inv1 g1097(.a(new_n1227_), .O(new_n1228_));
  nor2 g1098(.a(new_n1228_), .b(new_n1219_), .O(o_9_));
  inv1 g1099(.a(i_47_), .O(new_n1230_));
  nor2 g1100(.a(new_n393_), .b(new_n1230_), .O(new_n1231_));
  inv1 g1101(.a(new_n1231_), .O(new_n1232_));
  nor2 g1102(.a(new_n1232_), .b(new_n519_), .O(new_n1233_));
  inv1 g1103(.a(new_n1233_), .O(new_n1234_));
  nor2 g1104(.a(new_n1234_), .b(new_n935_), .O(o_62_));
  inv1 g1105(.a(i_56_), .O(new_n1236_));
  nor2 g1106(.a(new_n748_), .b(new_n1236_), .O(new_n1237_));
  inv1 g1107(.a(new_n1237_), .O(new_n1238_));
  nor2 g1108(.a(new_n1238_), .b(new_n935_), .O(o_63_));
  inv1 g1109(.a(i_53_), .O(new_n1240_));
  nor2 g1110(.a(new_n188_), .b(new_n1240_), .O(new_n1241_));
  inv1 g1111(.a(new_n1241_), .O(new_n1242_));
  nor2 g1112(.a(new_n1242_), .b(new_n827_), .O(new_n1243_));
  inv1 g1113(.a(new_n1243_), .O(new_n1244_));
  nor2 g1114(.a(new_n1244_), .b(new_n821_), .O(o_49_));
  inv1 g1115(.a(i_43_), .O(new_n1246_));
  nor2 g1116(.a(new_n1246_), .b(i_15_), .O(new_n1247_));
  inv1 g1117(.a(new_n1247_), .O(new_n1248_));
  nor2 g1118(.a(new_n1248_), .b(new_n411_), .O(o_7_));
  inv1 g1119(.a(i_30_), .O(new_n1250_));
  nor2 g1120(.a(new_n748_), .b(new_n1250_), .O(new_n1251_));
  inv1 g1121(.a(new_n1251_), .O(new_n1252_));
  nor2 g1122(.a(new_n1252_), .b(new_n755_), .O(new_n1253_));
  inv1 g1123(.a(new_n1253_), .O(new_n1254_));
  nor2 g1124(.a(new_n1254_), .b(new_n415_), .O(o_64_));
  inv1 g1125(.a(i_38_), .O(new_n1256_));
  nor2 g1126(.a(new_n155_), .b(new_n1256_), .O(new_n1257_));
  inv1 g1127(.a(new_n1257_), .O(new_n1258_));
  nor2 g1128(.a(new_n1258_), .b(new_n387_), .O(new_n1259_));
  inv1 g1129(.a(new_n1259_), .O(new_n1260_));
  nor2 g1130(.a(new_n1260_), .b(new_n623_), .O(new_n1261_));
  inv1 g1131(.a(new_n1261_), .O(new_n1262_));
  nor2 g1132(.a(new_n1262_), .b(new_n1091_), .O(new_n1263_));
  inv1 g1133(.a(new_n1263_), .O(new_n1264_));
  nor2 g1134(.a(new_n1215_), .b(new_n854_), .O(new_n1265_));
  inv1 g1135(.a(new_n1265_), .O(new_n1266_));
  nor2 g1136(.a(new_n1266_), .b(new_n1264_), .O(new_n1267_));
  inv1 g1137(.a(new_n1267_), .O(new_n1268_));
  nor2 g1138(.a(new_n1268_), .b(new_n335_), .O(o_8_));
  inv1 g1139(.a(i_40_), .O(new_n1270_));
  nor2 g1140(.a(new_n420_), .b(new_n1270_), .O(new_n1271_));
  inv1 g1141(.a(new_n1271_), .O(new_n1272_));
  nor2 g1142(.a(new_n1272_), .b(new_n713_), .O(o_59_));
  inv1 g1143(.a(i_14_), .O(new_n1274_));
  nor2 g1144(.a(i_15_), .b(new_n1274_), .O(new_n1275_));
  inv1 g1145(.a(new_n1275_), .O(new_n1276_));
  nor2 g1146(.a(new_n1276_), .b(new_n413_), .O(o_6_));
  nor2 g1147(.a(i_45_), .b(i_64_), .O(new_n1278_));
  inv1 g1148(.a(new_n1278_), .O(new_n1279_));
  inv1 g1149(.a(i_44_), .O(new_n1280_));
  nor2 g1150(.a(new_n1280_), .b(i_38_), .O(new_n1281_));
  inv1 g1151(.a(new_n1281_), .O(new_n1282_));
  nor2 g1152(.a(new_n1282_), .b(new_n1279_), .O(new_n1283_));
  inv1 g1153(.a(new_n1283_), .O(new_n1284_));
  nor2 g1154(.a(new_n1284_), .b(new_n547_), .O(new_n1285_));
  inv1 g1155(.a(new_n1285_), .O(new_n1286_));
  nor2 g1156(.a(new_n1286_), .b(new_n275_), .O(new_n1287_));
  inv1 g1157(.a(new_n1287_), .O(new_n1288_));
  nor2 g1158(.a(new_n1288_), .b(new_n561_), .O(new_n1289_));
  inv1 g1159(.a(new_n1289_), .O(new_n1290_));
  nor2 g1160(.a(new_n1215_), .b(new_n916_), .O(new_n1291_));
  inv1 g1161(.a(new_n1291_), .O(new_n1292_));
  nor2 g1162(.a(new_n1292_), .b(new_n1290_), .O(new_n1293_));
  inv1 g1163(.a(new_n1293_), .O(new_n1294_));
  nor2 g1164(.a(new_n1294_), .b(new_n335_), .O(o_3_));
  inv1 g1165(.a(i_15_), .O(new_n1296_));
  nor2 g1166(.a(new_n135_), .b(new_n1296_), .O(o_4_));
  buf  g1167(.a(i_29_), .O(o_5_));
endmodule


