// Benchmark "top" written by ABC on Wed Jan 17 21:32:51 2024

module top ( 
    i_89_, i_76_, i_63_, i_50_, i_75_, i_64_, i_78_, i_61_, i_99_, i_77_,
    i_62_, i_40_, i_72_, i_67_, i_71_, i_68_, i_74_, i_65_, i_30_, i_73_,
    i_66_, i_94_, i_81_, i_93_, i_82_, i_20_, i_92_, i_83_, i_69_, i_9_,
    i_91_, i_84_, i_98_, i_85_, i_10_, i_7_, i_97_, i_86_, i_79_, i_8_,
    i_96_, i_87_, i_5_, i_95_, i_88_, i_6_, i_27_, i_14_, i_3_, i_39_,
    i_28_, i_13_, i_4_, i_108_, i_25_, i_12_, i_1_, i_109_, i_26_, i_11_,
    i_2_, i_106_, i_90_, i_49_, i_23_, i_18_, i_116_, i_107_, i_24_, i_17_,
    i_0_, i_115_, i_104_, i_21_, i_16_, i_114_, i_105_, i_80_, i_59_,
    i_22_, i_15_, i_113_, i_102_, i_58_, i_45_, i_32_, i_112_, i_103_,
    i_57_, i_46_, i_31_, i_111_, i_100_, i_70_, i_56_, i_47_, i_34_,
    i_110_, i_101_, i_55_, i_48_, i_33_, i_19_, i_54_, i_41_, i_36_, i_60_,
    i_53_, i_42_, i_35_, i_52_, i_43_, i_38_, i_29_, i_51_, i_44_, i_37_,
    o_1_, o_80_, o_19_, o_2_, o_0_, o_70_, o_29_, o_60_, o_39_, o_38_,
    o_25_, o_12_, o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_,
    o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_,
    o_23_, o_18_, o_31_, o_24_, o_17_, o_69_, o_56_, o_43_, o_30_, o_55_,
    o_44_, o_58_, o_41_, o_79_, o_57_, o_42_, o_20_, o_52_, o_47_, o_51_,
    o_48_, o_54_, o_45_, o_10_, o_53_, o_46_, o_87_, o_74_, o_61_, o_9_,
    o_73_, o_62_, o_85_, o_72_, o_63_, o_49_, o_7_, o_86_, o_71_, o_64_,
    o_8_, o_83_, o_78_, o_65_, o_5_, o_84_, o_77_, o_66_, o_59_, o_6_,
    o_81_, o_76_, o_67_, o_3_, o_82_, o_75_, o_68_, o_4_  );
  input  i_89_, i_76_, i_63_, i_50_, i_75_, i_64_, i_78_, i_61_, i_99_,
    i_77_, i_62_, i_40_, i_72_, i_67_, i_71_, i_68_, i_74_, i_65_, i_30_,
    i_73_, i_66_, i_94_, i_81_, i_93_, i_82_, i_20_, i_92_, i_83_, i_69_,
    i_9_, i_91_, i_84_, i_98_, i_85_, i_10_, i_7_, i_97_, i_86_, i_79_,
    i_8_, i_96_, i_87_, i_5_, i_95_, i_88_, i_6_, i_27_, i_14_, i_3_,
    i_39_, i_28_, i_13_, i_4_, i_108_, i_25_, i_12_, i_1_, i_109_, i_26_,
    i_11_, i_2_, i_106_, i_90_, i_49_, i_23_, i_18_, i_116_, i_107_, i_24_,
    i_17_, i_0_, i_115_, i_104_, i_21_, i_16_, i_114_, i_105_, i_80_,
    i_59_, i_22_, i_15_, i_113_, i_102_, i_58_, i_45_, i_32_, i_112_,
    i_103_, i_57_, i_46_, i_31_, i_111_, i_100_, i_70_, i_56_, i_47_,
    i_34_, i_110_, i_101_, i_55_, i_48_, i_33_, i_19_, i_54_, i_41_, i_36_,
    i_60_, i_53_, i_42_, i_35_, i_52_, i_43_, i_38_, i_29_, i_51_, i_44_,
    i_37_;
  output o_1_, o_80_, o_19_, o_2_, o_0_, o_70_, o_29_, o_60_, o_39_, o_38_,
    o_25_, o_12_, o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_,
    o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_,
    o_23_, o_18_, o_31_, o_24_, o_17_, o_69_, o_56_, o_43_, o_30_, o_55_,
    o_44_, o_58_, o_41_, o_79_, o_57_, o_42_, o_20_, o_52_, o_47_, o_51_,
    o_48_, o_54_, o_45_, o_10_, o_53_, o_46_, o_87_, o_74_, o_61_, o_9_,
    o_73_, o_62_, o_85_, o_72_, o_63_, o_49_, o_7_, o_86_, o_71_, o_64_,
    o_8_, o_83_, o_78_, o_65_, o_5_, o_84_, o_77_, o_66_, o_59_, o_6_,
    o_81_, o_76_, o_67_, o_3_, o_82_, o_75_, o_68_, o_4_;
  wire new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n985_, new_n986_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1015_, new_n1016_, new_n1017_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1045_, new_n1046_,
    new_n1047_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_;
  nor2 g0000(.a(i_96_), .b(i_97_), .O(new_n206_));
  inv1 g0001(.a(new_n206_), .O(new_n207_));
  nor2 g0002(.a(i_100_), .b(i_95_), .O(new_n208_));
  inv1 g0003(.a(new_n208_), .O(new_n209_));
  nor2 g0004(.a(new_n209_), .b(new_n207_), .O(new_n210_));
  inv1 g0005(.a(new_n210_), .O(new_n211_));
  nor2 g0006(.a(i_94_), .b(i_99_), .O(new_n212_));
  inv1 g0007(.a(new_n212_), .O(new_n213_));
  nor2 g0008(.a(i_98_), .b(i_93_), .O(new_n214_));
  inv1 g0009(.a(new_n214_), .O(new_n215_));
  nor2 g0010(.a(new_n215_), .b(new_n213_), .O(new_n216_));
  inv1 g0011(.a(new_n216_), .O(new_n217_));
  nor2 g0012(.a(new_n217_), .b(new_n211_), .O(new_n218_));
  inv1 g0013(.a(new_n218_), .O(o_1_));
  inv1 g0014(.a(i_3_), .O(new_n220_));
  inv1 g0015(.a(i_30_), .O(new_n221_));
  inv1 g0016(.a(i_29_), .O(new_n222_));
  nor2 g0017(.a(new_n222_), .b(new_n221_), .O(new_n223_));
  inv1 g0018(.a(new_n223_), .O(new_n224_));
  nor2 g0019(.a(new_n224_), .b(new_n220_), .O(new_n225_));
  inv1 g0020(.a(new_n225_), .O(new_n226_));
  inv1 g0021(.a(i_4_), .O(new_n227_));
  inv1 g0022(.a(i_32_), .O(new_n228_));
  inv1 g0023(.a(i_31_), .O(new_n229_));
  nor2 g0024(.a(new_n229_), .b(new_n228_), .O(new_n230_));
  inv1 g0025(.a(new_n230_), .O(new_n231_));
  nor2 g0026(.a(new_n231_), .b(new_n227_), .O(new_n232_));
  inv1 g0027(.a(new_n232_), .O(new_n233_));
  nor2 g0028(.a(new_n233_), .b(new_n226_), .O(new_n234_));
  inv1 g0029(.a(new_n234_), .O(new_n235_));
  nor2 g0030(.a(new_n235_), .b(i_33_), .O(new_n236_));
  inv1 g0031(.a(new_n236_), .O(new_n237_));
  inv1 g0032(.a(i_108_), .O(new_n238_));
  inv1 g0033(.a(i_107_), .O(new_n239_));
  nor2 g0034(.a(new_n239_), .b(new_n238_), .O(new_n240_));
  inv1 g0035(.a(new_n240_), .O(new_n241_));
  inv1 g0036(.a(i_106_), .O(new_n242_));
  inv1 g0037(.a(i_105_), .O(new_n243_));
  nor2 g0038(.a(new_n243_), .b(new_n242_), .O(new_n244_));
  inv1 g0039(.a(new_n244_), .O(new_n245_));
  nor2 g0040(.a(new_n245_), .b(new_n241_), .O(new_n246_));
  inv1 g0041(.a(new_n246_), .O(new_n247_));
  inv1 g0042(.a(i_104_), .O(new_n248_));
  inv1 g0043(.a(i_101_), .O(new_n249_));
  inv1 g0044(.a(i_102_), .O(new_n250_));
  inv1 g0045(.a(i_103_), .O(new_n251_));
  nor2 g0046(.a(new_n251_), .b(new_n250_), .O(new_n252_));
  inv1 g0047(.a(new_n252_), .O(new_n253_));
  nor2 g0048(.a(new_n253_), .b(new_n249_), .O(new_n254_));
  inv1 g0049(.a(new_n254_), .O(new_n255_));
  nor2 g0050(.a(new_n255_), .b(new_n248_), .O(new_n256_));
  inv1 g0051(.a(new_n256_), .O(new_n257_));
  nor2 g0052(.a(new_n257_), .b(new_n247_), .O(new_n258_));
  inv1 g0053(.a(new_n258_), .O(new_n259_));
  nor2 g0054(.a(new_n259_), .b(i_109_), .O(new_n260_));
  inv1 g0055(.a(new_n260_), .O(new_n261_));
  nor2 g0056(.a(new_n261_), .b(new_n237_), .O(new_n262_));
  inv1 g0057(.a(i_6_), .O(new_n263_));
  nor2 g0058(.a(new_n227_), .b(new_n263_), .O(new_n264_));
  inv1 g0059(.a(new_n264_), .O(new_n265_));
  nor2 g0060(.a(new_n226_), .b(new_n229_), .O(new_n266_));
  inv1 g0061(.a(new_n266_), .O(new_n267_));
  nor2 g0062(.a(new_n267_), .b(new_n265_), .O(new_n268_));
  inv1 g0063(.a(new_n268_), .O(new_n269_));
  inv1 g0064(.a(i_114_), .O(new_n270_));
  inv1 g0065(.a(i_110_), .O(new_n271_));
  nor2 g0066(.a(new_n271_), .b(new_n270_), .O(new_n272_));
  inv1 g0067(.a(new_n272_), .O(new_n273_));
  inv1 g0068(.a(i_113_), .O(new_n274_));
  inv1 g0069(.a(i_112_), .O(new_n275_));
  inv1 g0070(.a(i_111_), .O(new_n276_));
  nor2 g0071(.a(new_n276_), .b(new_n275_), .O(new_n277_));
  inv1 g0072(.a(new_n277_), .O(new_n278_));
  inv1 g0073(.a(i_116_), .O(new_n279_));
  inv1 g0074(.a(i_115_), .O(new_n280_));
  nor2 g0075(.a(new_n280_), .b(new_n279_), .O(new_n281_));
  inv1 g0076(.a(new_n281_), .O(new_n282_));
  nor2 g0077(.a(new_n282_), .b(new_n278_), .O(new_n283_));
  inv1 g0078(.a(new_n283_), .O(new_n284_));
  nor2 g0079(.a(new_n284_), .b(new_n274_), .O(new_n285_));
  inv1 g0080(.a(new_n285_), .O(new_n286_));
  nor2 g0081(.a(new_n286_), .b(new_n273_), .O(new_n287_));
  nor2 g0082(.a(new_n253_), .b(new_n248_), .O(new_n288_));
  inv1 g0083(.a(new_n288_), .O(new_n289_));
  nor2 g0084(.a(new_n289_), .b(new_n247_), .O(new_n290_));
  inv1 g0085(.a(new_n290_), .O(new_n291_));
  nor2 g0086(.a(i_33_), .b(new_n228_), .O(new_n292_));
  inv1 g0087(.a(new_n292_), .O(new_n293_));
  nor2 g0088(.a(new_n293_), .b(new_n249_), .O(new_n294_));
  inv1 g0089(.a(new_n294_), .O(new_n295_));
  nor2 g0090(.a(new_n295_), .b(new_n291_), .O(new_n296_));
  inv1 g0091(.a(new_n296_), .O(new_n297_));
  nor2 g0092(.a(new_n297_), .b(new_n287_), .O(new_n298_));
  inv1 g0093(.a(new_n298_), .O(new_n299_));
  nor2 g0094(.a(new_n299_), .b(new_n269_), .O(new_n300_));
  inv1 g0095(.a(i_109_), .O(new_n301_));
  nor2 g0096(.a(new_n271_), .b(new_n301_), .O(new_n302_));
  inv1 g0097(.a(new_n302_), .O(new_n303_));
  nor2 g0098(.a(new_n303_), .b(new_n291_), .O(new_n304_));
  inv1 g0099(.a(new_n304_), .O(new_n305_));
  nor2 g0100(.a(new_n284_), .b(new_n249_), .O(new_n306_));
  inv1 g0101(.a(new_n306_), .O(new_n307_));
  nor2 g0102(.a(new_n307_), .b(new_n305_), .O(new_n308_));
  inv1 g0103(.a(new_n308_), .O(new_n309_));
  nor2 g0104(.a(new_n227_), .b(i_6_), .O(new_n310_));
  inv1 g0105(.a(new_n310_), .O(new_n311_));
  nor2 g0106(.a(new_n311_), .b(new_n274_), .O(new_n312_));
  inv1 g0107(.a(new_n312_), .O(new_n313_));
  nor2 g0108(.a(new_n313_), .b(new_n270_), .O(new_n314_));
  inv1 g0109(.a(new_n314_), .O(new_n315_));
  nor2 g0110(.a(new_n315_), .b(new_n309_), .O(new_n316_));
  nor2 g0111(.a(new_n316_), .b(new_n300_), .O(new_n317_));
  inv1 g0112(.a(new_n317_), .O(new_n318_));
  nor2 g0113(.a(new_n318_), .b(new_n262_), .O(new_n319_));
  inv1 g0114(.a(new_n319_), .O(new_n320_));
  inv1 g0115(.a(i_5_), .O(new_n321_));
  nor2 g0116(.a(new_n311_), .b(new_n321_), .O(new_n322_));
  inv1 g0117(.a(new_n322_), .O(new_n323_));
  nor2 g0118(.a(new_n323_), .b(new_n258_), .O(new_n324_));
  nor2 g0119(.a(new_n311_), .b(new_n236_), .O(new_n325_));
  nor2 g0120(.a(new_n325_), .b(new_n324_), .O(new_n326_));
  nor2 g0121(.a(new_n326_), .b(new_n301_), .O(new_n327_));
  nor2 g0122(.a(new_n231_), .b(i_33_), .O(new_n328_));
  inv1 g0123(.a(new_n328_), .O(new_n329_));
  nor2 g0124(.a(new_n329_), .b(new_n226_), .O(new_n330_));
  inv1 g0125(.a(new_n330_), .O(new_n331_));
  nor2 g0126(.a(new_n331_), .b(i_5_), .O(new_n332_));
  inv1 g0127(.a(new_n332_), .O(new_n333_));
  nor2 g0128(.a(new_n333_), .b(new_n265_), .O(new_n334_));
  inv1 g0129(.a(new_n334_), .O(new_n335_));
  inv1 g0130(.a(new_n287_), .O(new_n336_));
  nor2 g0131(.a(new_n336_), .b(new_n259_), .O(new_n337_));
  nor2 g0132(.a(new_n337_), .b(new_n335_), .O(new_n338_));
  nor2 g0133(.a(new_n237_), .b(i_5_), .O(new_n339_));
  inv1 g0134(.a(new_n339_), .O(new_n340_));
  nor2 g0135(.a(new_n340_), .b(i_109_), .O(new_n341_));
  nor2 g0136(.a(new_n341_), .b(new_n338_), .O(new_n342_));
  inv1 g0137(.a(new_n342_), .O(new_n343_));
  nor2 g0138(.a(new_n343_), .b(new_n327_), .O(new_n344_));
  inv1 g0139(.a(new_n344_), .O(new_n345_));
  nor2 g0140(.a(new_n345_), .b(new_n320_), .O(new_n346_));
  inv1 g0141(.a(new_n346_), .O(o_80_));
  inv1 g0142(.a(i_1_), .O(new_n348_));
  nor2 g0143(.a(new_n348_), .b(new_n227_), .O(new_n349_));
  inv1 g0144(.a(new_n349_), .O(new_n350_));
  nor2 g0145(.a(new_n350_), .b(i_0_), .O(new_n351_));
  inv1 g0146(.a(new_n351_), .O(new_n352_));
  nor2 g0147(.a(new_n352_), .b(i_28_), .O(new_n353_));
  nor2 g0148(.a(new_n351_), .b(i_36_), .O(new_n354_));
  nor2 g0149(.a(new_n354_), .b(new_n353_), .O(o_2_));
  nor2 g0150(.a(new_n329_), .b(new_n224_), .O(new_n356_));
  inv1 g0151(.a(new_n356_), .O(new_n357_));
  nor2 g0152(.a(new_n348_), .b(i_28_), .O(new_n358_));
  inv1 g0153(.a(new_n358_), .O(new_n359_));
  nor2 g0154(.a(i_26_), .b(i_27_), .O(new_n360_));
  inv1 g0155(.a(new_n360_), .O(new_n361_));
  nor2 g0156(.a(new_n361_), .b(new_n359_), .O(new_n362_));
  inv1 g0157(.a(new_n362_), .O(new_n363_));
  nor2 g0158(.a(new_n363_), .b(i_25_), .O(new_n364_));
  nor2 g0159(.a(new_n364_), .b(new_n357_), .O(new_n365_));
  inv1 g0160(.a(new_n365_), .O(new_n366_));
  nor2 g0161(.a(new_n366_), .b(new_n227_), .O(new_n367_));
  nor2 g0162(.a(i_24_), .b(i_23_), .O(new_n368_));
  inv1 g0163(.a(new_n368_), .O(new_n369_));
  nor2 g0164(.a(new_n369_), .b(new_n227_), .O(new_n370_));
  inv1 g0165(.a(new_n370_), .O(new_n371_));
  nor2 g0166(.a(new_n371_), .b(new_n357_), .O(new_n372_));
  inv1 g0167(.a(i_0_), .O(new_n373_));
  nor2 g0168(.a(new_n373_), .b(new_n227_), .O(new_n374_));
  inv1 g0169(.a(new_n374_), .O(new_n375_));
  inv1 g0170(.a(i_23_), .O(new_n376_));
  nor2 g0171(.a(i_24_), .b(new_n376_), .O(new_n377_));
  nor2 g0172(.a(i_0_), .b(i_23_), .O(new_n378_));
  nor2 g0173(.a(new_n378_), .b(new_n377_), .O(new_n379_));
  inv1 g0174(.a(new_n379_), .O(new_n380_));
  nor2 g0175(.a(new_n380_), .b(new_n357_), .O(new_n381_));
  inv1 g0176(.a(new_n381_), .O(new_n382_));
  nor2 g0177(.a(new_n382_), .b(new_n375_), .O(new_n383_));
  nor2 g0178(.a(new_n383_), .b(new_n372_), .O(new_n384_));
  inv1 g0179(.a(new_n384_), .O(new_n385_));
  nor2 g0180(.a(new_n385_), .b(new_n367_), .O(new_n386_));
  nor2 g0181(.a(i_13_), .b(i_91_), .O(new_n387_));
  inv1 g0182(.a(i_91_), .O(new_n388_));
  inv1 g0183(.a(i_13_), .O(new_n389_));
  nor2 g0184(.a(new_n389_), .b(new_n388_), .O(new_n390_));
  nor2 g0185(.a(new_n390_), .b(new_n387_), .O(new_n391_));
  inv1 g0186(.a(new_n391_), .O(new_n392_));
  nor2 g0187(.a(new_n392_), .b(i_83_), .O(new_n393_));
  inv1 g0188(.a(new_n393_), .O(new_n394_));
  nor2 g0189(.a(new_n394_), .b(new_n386_), .O(new_n395_));
  nor2 g0190(.a(new_n231_), .b(new_n224_), .O(new_n396_));
  inv1 g0191(.a(new_n396_), .O(new_n397_));
  inv1 g0192(.a(i_24_), .O(new_n398_));
  inv1 g0193(.a(new_n353_), .O(new_n399_));
  nor2 g0194(.a(i_25_), .b(i_27_), .O(new_n400_));
  inv1 g0195(.a(new_n400_), .O(new_n401_));
  nor2 g0196(.a(new_n401_), .b(i_26_), .O(new_n402_));
  inv1 g0197(.a(new_n402_), .O(new_n403_));
  nor2 g0198(.a(new_n403_), .b(new_n399_), .O(new_n404_));
  inv1 g0199(.a(new_n404_), .O(new_n405_));
  nor2 g0200(.a(new_n405_), .b(new_n398_), .O(new_n406_));
  inv1 g0201(.a(new_n406_), .O(new_n407_));
  nor2 g0202(.a(new_n407_), .b(new_n397_), .O(new_n408_));
  inv1 g0203(.a(new_n408_), .O(new_n409_));
  nor2 g0204(.a(new_n391_), .b(i_23_), .O(new_n410_));
  nor2 g0205(.a(new_n389_), .b(i_83_), .O(new_n411_));
  nor2 g0206(.a(new_n411_), .b(new_n376_), .O(new_n412_));
  nor2 g0207(.a(i_33_), .b(i_21_), .O(new_n413_));
  inv1 g0208(.a(new_n413_), .O(new_n414_));
  nor2 g0209(.a(new_n414_), .b(new_n412_), .O(new_n415_));
  inv1 g0210(.a(new_n415_), .O(new_n416_));
  nor2 g0211(.a(new_n416_), .b(new_n410_), .O(new_n417_));
  inv1 g0212(.a(new_n417_), .O(new_n418_));
  nor2 g0213(.a(new_n418_), .b(new_n409_), .O(new_n419_));
  inv1 g0214(.a(i_99_), .O(new_n420_));
  inv1 g0215(.a(new_n377_), .O(new_n421_));
  nor2 g0216(.a(new_n421_), .b(i_25_), .O(new_n422_));
  inv1 g0217(.a(new_n422_), .O(new_n423_));
  nor2 g0218(.a(new_n363_), .b(i_0_), .O(new_n424_));
  inv1 g0219(.a(new_n424_), .O(new_n425_));
  nor2 g0220(.a(new_n425_), .b(new_n423_), .O(new_n426_));
  nor2 g0221(.a(new_n426_), .b(new_n227_), .O(new_n427_));
  inv1 g0222(.a(new_n427_), .O(new_n428_));
  nor2 g0223(.a(new_n428_), .b(new_n420_), .O(new_n429_));
  inv1 g0224(.a(i_21_), .O(new_n430_));
  nor2 g0225(.a(new_n421_), .b(new_n430_), .O(new_n431_));
  nor2 g0226(.a(new_n430_), .b(new_n376_), .O(new_n432_));
  inv1 g0227(.a(new_n432_), .O(new_n433_));
  nor2 g0228(.a(i_13_), .b(i_83_), .O(new_n434_));
  inv1 g0229(.a(new_n434_), .O(new_n435_));
  nor2 g0230(.a(new_n435_), .b(new_n433_), .O(new_n436_));
  inv1 g0231(.a(new_n436_), .O(new_n437_));
  nor2 g0232(.a(new_n437_), .b(new_n357_), .O(new_n438_));
  nor2 g0233(.a(new_n438_), .b(new_n431_), .O(new_n439_));
  nor2 g0234(.a(new_n439_), .b(new_n405_), .O(new_n440_));
  nor2 g0235(.a(new_n440_), .b(new_n429_), .O(new_n441_));
  inv1 g0236(.a(new_n441_), .O(new_n442_));
  nor2 g0237(.a(new_n442_), .b(new_n419_), .O(new_n443_));
  inv1 g0238(.a(new_n443_), .O(new_n444_));
  nor2 g0239(.a(new_n444_), .b(new_n395_), .O(new_n445_));
  inv1 g0240(.a(new_n445_), .O(o_70_));
  inv1 g0241(.a(i_89_), .O(new_n448_));
  nor2 g0242(.a(new_n407_), .b(new_n376_), .O(new_n449_));
  nor2 g0243(.a(new_n449_), .b(new_n227_), .O(new_n450_));
  inv1 g0244(.a(new_n450_), .O(new_n451_));
  nor2 g0245(.a(new_n451_), .b(new_n448_), .O(new_n452_));
  inv1 g0246(.a(i_19_), .O(new_n453_));
  inv1 g0247(.a(new_n449_), .O(new_n454_));
  nor2 g0248(.a(new_n454_), .b(new_n453_), .O(new_n455_));
  nor2 g0249(.a(new_n455_), .b(new_n452_), .O(new_n456_));
  inv1 g0250(.a(new_n456_), .O(o_60_));
  inv1 g0251(.a(i_68_), .O(new_n458_));
  nor2 g0252(.a(new_n369_), .b(i_25_), .O(new_n459_));
  inv1 g0253(.a(new_n459_), .O(new_n460_));
  inv1 g0254(.a(i_26_), .O(new_n461_));
  nor2 g0255(.a(new_n461_), .b(i_27_), .O(new_n462_));
  inv1 g0256(.a(new_n462_), .O(new_n463_));
  nor2 g0257(.a(new_n463_), .b(new_n359_), .O(new_n464_));
  inv1 g0258(.a(new_n464_), .O(new_n465_));
  nor2 g0259(.a(new_n465_), .b(new_n460_), .O(new_n466_));
  nor2 g0260(.a(new_n466_), .b(new_n311_), .O(new_n467_));
  nor2 g0261(.a(new_n460_), .b(new_n375_), .O(new_n468_));
  inv1 g0262(.a(new_n468_), .O(new_n469_));
  nor2 g0263(.a(new_n469_), .b(new_n465_), .O(new_n470_));
  nor2 g0264(.a(new_n470_), .b(new_n467_), .O(new_n471_));
  nor2 g0265(.a(new_n471_), .b(new_n458_), .O(new_n472_));
  nor2 g0266(.a(new_n466_), .b(new_n265_), .O(new_n473_));
  inv1 g0267(.a(new_n473_), .O(new_n474_));
  nor2 g0268(.a(new_n474_), .b(new_n238_), .O(new_n475_));
  inv1 g0269(.a(i_22_), .O(new_n476_));
  nor2 g0270(.a(new_n369_), .b(new_n476_), .O(new_n477_));
  inv1 g0271(.a(new_n477_), .O(new_n478_));
  nor2 g0272(.a(new_n401_), .b(new_n461_), .O(new_n479_));
  inv1 g0273(.a(new_n479_), .O(new_n480_));
  nor2 g0274(.a(new_n480_), .b(new_n399_), .O(new_n481_));
  inv1 g0275(.a(new_n481_), .O(new_n482_));
  nor2 g0276(.a(new_n482_), .b(new_n478_), .O(new_n483_));
  nor2 g0277(.a(new_n483_), .b(new_n475_), .O(new_n484_));
  inv1 g0278(.a(new_n484_), .O(new_n485_));
  nor2 g0279(.a(new_n485_), .b(new_n472_), .O(new_n486_));
  inv1 g0280(.a(new_n486_), .O(o_39_));
  inv1 g0281(.a(i_67_), .O(new_n488_));
  nor2 g0282(.a(new_n471_), .b(new_n488_), .O(new_n489_));
  nor2 g0283(.a(new_n474_), .b(new_n239_), .O(new_n490_));
  nor2 g0284(.a(new_n369_), .b(new_n430_), .O(new_n491_));
  inv1 g0285(.a(new_n491_), .O(new_n492_));
  nor2 g0286(.a(new_n492_), .b(new_n482_), .O(new_n493_));
  nor2 g0287(.a(new_n493_), .b(new_n490_), .O(new_n494_));
  inv1 g0288(.a(new_n494_), .O(new_n495_));
  nor2 g0289(.a(new_n495_), .b(new_n489_), .O(new_n496_));
  inv1 g0290(.a(new_n496_), .O(o_38_));
  inv1 g0291(.a(i_57_), .O(new_n498_));
  inv1 g0292(.a(i_25_), .O(new_n499_));
  nor2 g0293(.a(new_n369_), .b(new_n499_), .O(new_n500_));
  inv1 g0294(.a(new_n500_), .O(new_n501_));
  nor2 g0295(.a(new_n501_), .b(new_n425_), .O(new_n502_));
  nor2 g0296(.a(new_n502_), .b(new_n227_), .O(new_n503_));
  inv1 g0297(.a(new_n503_), .O(new_n504_));
  nor2 g0298(.a(new_n504_), .b(new_n498_), .O(new_n505_));
  nor2 g0299(.a(new_n369_), .b(new_n453_), .O(new_n506_));
  inv1 g0300(.a(new_n506_), .O(new_n507_));
  nor2 g0301(.a(new_n361_), .b(new_n499_), .O(new_n508_));
  inv1 g0302(.a(new_n508_), .O(new_n509_));
  nor2 g0303(.a(new_n509_), .b(new_n399_), .O(new_n510_));
  inv1 g0304(.a(new_n510_), .O(new_n511_));
  nor2 g0305(.a(new_n511_), .b(new_n507_), .O(new_n512_));
  nor2 g0306(.a(new_n512_), .b(new_n505_), .O(new_n513_));
  inv1 g0307(.a(new_n513_), .O(o_25_));
  inv1 g0308(.a(i_27_), .O(new_n515_));
  nor2 g0309(.a(i_25_), .b(new_n515_), .O(new_n516_));
  inv1 g0310(.a(new_n516_), .O(new_n517_));
  nor2 g0311(.a(new_n517_), .b(i_26_), .O(new_n518_));
  inv1 g0312(.a(new_n518_), .O(new_n519_));
  inv1 g0313(.a(i_16_), .O(new_n520_));
  nor2 g0314(.a(new_n369_), .b(new_n520_), .O(new_n521_));
  inv1 g0315(.a(new_n521_), .O(new_n522_));
  nor2 g0316(.a(new_n522_), .b(new_n399_), .O(new_n523_));
  inv1 g0317(.a(new_n523_), .O(new_n524_));
  nor2 g0318(.a(new_n524_), .b(new_n519_), .O(new_n525_));
  inv1 g0319(.a(i_46_), .O(new_n526_));
  nor2 g0320(.a(i_26_), .b(new_n515_), .O(new_n527_));
  inv1 g0321(.a(new_n527_), .O(new_n528_));
  nor2 g0322(.a(new_n528_), .b(new_n359_), .O(new_n529_));
  inv1 g0323(.a(new_n529_), .O(new_n530_));
  nor2 g0324(.a(new_n460_), .b(i_0_), .O(new_n531_));
  inv1 g0325(.a(new_n531_), .O(new_n532_));
  nor2 g0326(.a(new_n532_), .b(new_n530_), .O(new_n533_));
  nor2 g0327(.a(new_n533_), .b(new_n227_), .O(new_n534_));
  inv1 g0328(.a(new_n534_), .O(new_n535_));
  nor2 g0329(.a(new_n535_), .b(new_n526_), .O(new_n536_));
  nor2 g0330(.a(new_n536_), .b(new_n525_), .O(new_n537_));
  inv1 g0331(.a(new_n537_), .O(o_12_));
  inv1 g0332(.a(i_66_), .O(new_n539_));
  nor2 g0333(.a(new_n471_), .b(new_n539_), .O(new_n540_));
  inv1 g0334(.a(i_20_), .O(new_n541_));
  nor2 g0335(.a(new_n369_), .b(new_n541_), .O(new_n542_));
  inv1 g0336(.a(new_n542_), .O(new_n543_));
  nor2 g0337(.a(new_n543_), .b(new_n482_), .O(new_n544_));
  nor2 g0338(.a(new_n474_), .b(new_n242_), .O(new_n545_));
  nor2 g0339(.a(new_n545_), .b(new_n544_), .O(new_n546_));
  inv1 g0340(.a(new_n546_), .O(new_n547_));
  nor2 g0341(.a(new_n547_), .b(new_n540_), .O(new_n548_));
  inv1 g0342(.a(new_n548_), .O(o_37_));
  nor2 g0343(.a(new_n543_), .b(new_n511_), .O(new_n550_));
  inv1 g0344(.a(i_58_), .O(new_n551_));
  nor2 g0345(.a(new_n504_), .b(new_n551_), .O(new_n552_));
  nor2 g0346(.a(new_n552_), .b(new_n550_), .O(new_n553_));
  inv1 g0347(.a(new_n553_), .O(o_26_));
  inv1 g0348(.a(i_45_), .O(new_n555_));
  nor2 g0349(.a(new_n535_), .b(new_n555_), .O(new_n556_));
  inv1 g0350(.a(i_15_), .O(new_n557_));
  nor2 g0351(.a(new_n369_), .b(new_n557_), .O(new_n558_));
  inv1 g0352(.a(new_n558_), .O(new_n559_));
  nor2 g0353(.a(new_n559_), .b(new_n399_), .O(new_n560_));
  inv1 g0354(.a(new_n560_), .O(new_n561_));
  nor2 g0355(.a(new_n561_), .b(new_n519_), .O(new_n562_));
  nor2 g0356(.a(new_n562_), .b(new_n556_), .O(new_n563_));
  inv1 g0357(.a(new_n563_), .O(o_11_));
  inv1 g0358(.a(i_79_), .O(new_n565_));
  nor2 g0359(.a(new_n398_), .b(i_25_), .O(new_n566_));
  inv1 g0360(.a(new_n566_), .O(new_n567_));
  nor2 g0361(.a(new_n567_), .b(i_23_), .O(new_n568_));
  inv1 g0362(.a(new_n568_), .O(new_n569_));
  nor2 g0363(.a(new_n569_), .b(new_n425_), .O(new_n570_));
  nor2 g0364(.a(new_n570_), .b(new_n565_), .O(new_n571_));
  inv1 g0365(.a(i_17_), .O(new_n572_));
  inv1 g0366(.a(new_n570_), .O(new_n573_));
  nor2 g0367(.a(new_n573_), .b(new_n572_), .O(new_n574_));
  nor2 g0368(.a(new_n574_), .b(new_n227_), .O(new_n575_));
  inv1 g0369(.a(new_n575_), .O(new_n576_));
  nor2 g0370(.a(new_n576_), .b(new_n571_), .O(new_n577_));
  inv1 g0371(.a(new_n577_), .O(o_50_));
  inv1 g0372(.a(i_65_), .O(new_n579_));
  nor2 g0373(.a(new_n471_), .b(new_n579_), .O(new_n580_));
  nor2 g0374(.a(new_n507_), .b(new_n482_), .O(new_n581_));
  nor2 g0375(.a(new_n474_), .b(new_n243_), .O(new_n582_));
  nor2 g0376(.a(new_n582_), .b(new_n581_), .O(new_n583_));
  inv1 g0377(.a(new_n583_), .O(new_n584_));
  nor2 g0378(.a(new_n584_), .b(new_n580_), .O(new_n585_));
  inv1 g0379(.a(new_n585_), .O(o_36_));
  inv1 g0380(.a(i_35_), .O(new_n587_));
  nor2 g0381(.a(new_n587_), .b(new_n227_), .O(o_27_));
  inv1 g0382(.a(i_48_), .O(new_n589_));
  nor2 g0383(.a(new_n535_), .b(new_n589_), .O(new_n590_));
  inv1 g0384(.a(i_18_), .O(new_n591_));
  nor2 g0385(.a(new_n369_), .b(new_n591_), .O(new_n592_));
  inv1 g0386(.a(new_n592_), .O(new_n593_));
  nor2 g0387(.a(new_n593_), .b(new_n399_), .O(new_n594_));
  inv1 g0388(.a(new_n594_), .O(new_n595_));
  nor2 g0389(.a(new_n595_), .b(new_n519_), .O(new_n596_));
  nor2 g0390(.a(new_n596_), .b(new_n590_), .O(new_n597_));
  inv1 g0391(.a(new_n597_), .O(o_14_));
  inv1 g0392(.a(i_64_), .O(new_n599_));
  nor2 g0393(.a(new_n471_), .b(new_n599_), .O(new_n600_));
  nor2 g0394(.a(new_n595_), .b(new_n480_), .O(new_n601_));
  nor2 g0395(.a(new_n474_), .b(new_n248_), .O(new_n602_));
  nor2 g0396(.a(new_n602_), .b(new_n601_), .O(new_n603_));
  inv1 g0397(.a(new_n603_), .O(new_n604_));
  nor2 g0398(.a(new_n604_), .b(new_n600_), .O(new_n605_));
  inv1 g0399(.a(new_n605_), .O(o_35_));
  inv1 g0400(.a(i_34_), .O(new_n607_));
  nor2 g0401(.a(new_n607_), .b(new_n227_), .O(o_28_));
  inv1 g0402(.a(i_47_), .O(new_n609_));
  nor2 g0403(.a(new_n535_), .b(new_n609_), .O(new_n610_));
  nor2 g0404(.a(new_n369_), .b(new_n572_), .O(new_n611_));
  inv1 g0405(.a(new_n611_), .O(new_n612_));
  nor2 g0406(.a(new_n612_), .b(new_n399_), .O(new_n613_));
  inv1 g0407(.a(new_n613_), .O(new_n614_));
  nor2 g0408(.a(new_n614_), .b(new_n519_), .O(new_n615_));
  nor2 g0409(.a(new_n615_), .b(new_n610_), .O(new_n616_));
  inv1 g0410(.a(new_n616_), .O(o_13_));
  inv1 g0411(.a(i_63_), .O(new_n618_));
  nor2 g0412(.a(new_n471_), .b(new_n618_), .O(new_n619_));
  nor2 g0413(.a(new_n614_), .b(new_n480_), .O(new_n620_));
  nor2 g0414(.a(new_n474_), .b(new_n251_), .O(new_n621_));
  nor2 g0415(.a(new_n621_), .b(new_n620_), .O(new_n622_));
  inv1 g0416(.a(new_n622_), .O(new_n623_));
  nor2 g0417(.a(new_n623_), .b(new_n619_), .O(new_n624_));
  inv1 g0418(.a(new_n624_), .O(o_34_));
  inv1 g0419(.a(i_53_), .O(new_n626_));
  nor2 g0420(.a(new_n504_), .b(new_n626_), .O(new_n627_));
  nor2 g0421(.a(new_n561_), .b(new_n509_), .O(new_n628_));
  nor2 g0422(.a(new_n628_), .b(new_n627_), .O(new_n629_));
  inv1 g0423(.a(new_n629_), .O(o_21_));
  inv1 g0424(.a(i_50_), .O(new_n631_));
  nor2 g0425(.a(new_n535_), .b(new_n631_), .O(new_n632_));
  nor2 g0426(.a(new_n519_), .b(new_n399_), .O(new_n633_));
  inv1 g0427(.a(new_n633_), .O(new_n634_));
  nor2 g0428(.a(new_n634_), .b(new_n543_), .O(new_n635_));
  nor2 g0429(.a(new_n635_), .b(new_n632_), .O(new_n636_));
  inv1 g0430(.a(new_n636_), .O(o_16_));
  inv1 g0431(.a(i_69_), .O(new_n638_));
  nor2 g0432(.a(new_n465_), .b(new_n423_), .O(new_n639_));
  nor2 g0433(.a(new_n639_), .b(new_n311_), .O(new_n640_));
  inv1 g0434(.a(new_n639_), .O(new_n641_));
  nor2 g0435(.a(new_n641_), .b(new_n375_), .O(new_n642_));
  nor2 g0436(.a(new_n642_), .b(new_n640_), .O(new_n643_));
  nor2 g0437(.a(new_n643_), .b(new_n638_), .O(new_n644_));
  nor2 g0438(.a(new_n639_), .b(new_n265_), .O(new_n645_));
  inv1 g0439(.a(new_n645_), .O(new_n646_));
  nor2 g0440(.a(new_n646_), .b(new_n301_), .O(new_n647_));
  nor2 g0441(.a(new_n421_), .b(new_n557_), .O(new_n648_));
  inv1 g0442(.a(new_n648_), .O(new_n649_));
  nor2 g0443(.a(new_n649_), .b(new_n482_), .O(new_n650_));
  nor2 g0444(.a(new_n650_), .b(new_n647_), .O(new_n651_));
  inv1 g0445(.a(new_n651_), .O(new_n652_));
  nor2 g0446(.a(new_n652_), .b(new_n644_), .O(new_n653_));
  inv1 g0447(.a(new_n653_), .O(o_40_));
  inv1 g0448(.a(i_62_), .O(new_n655_));
  nor2 g0449(.a(new_n471_), .b(new_n655_), .O(new_n656_));
  nor2 g0450(.a(new_n524_), .b(new_n480_), .O(new_n657_));
  nor2 g0451(.a(new_n474_), .b(new_n250_), .O(new_n658_));
  nor2 g0452(.a(new_n658_), .b(new_n657_), .O(new_n659_));
  inv1 g0453(.a(new_n659_), .O(new_n660_));
  nor2 g0454(.a(new_n660_), .b(new_n656_), .O(new_n661_));
  inv1 g0455(.a(new_n661_), .O(o_33_));
  inv1 g0456(.a(i_54_), .O(new_n663_));
  nor2 g0457(.a(new_n504_), .b(new_n663_), .O(new_n664_));
  nor2 g0458(.a(new_n524_), .b(new_n509_), .O(new_n665_));
  nor2 g0459(.a(new_n665_), .b(new_n664_), .O(new_n666_));
  inv1 g0460(.a(new_n666_), .O(o_22_));
  inv1 g0461(.a(i_49_), .O(new_n668_));
  nor2 g0462(.a(new_n535_), .b(new_n668_), .O(new_n669_));
  nor2 g0463(.a(new_n634_), .b(new_n507_), .O(new_n670_));
  nor2 g0464(.a(new_n670_), .b(new_n669_), .O(new_n671_));
  inv1 g0465(.a(new_n671_), .O(o_15_));
  inv1 g0466(.a(i_61_), .O(new_n673_));
  nor2 g0467(.a(new_n471_), .b(new_n673_), .O(new_n674_));
  nor2 g0468(.a(new_n474_), .b(new_n249_), .O(new_n675_));
  nor2 g0469(.a(new_n561_), .b(new_n480_), .O(new_n676_));
  nor2 g0470(.a(new_n676_), .b(new_n675_), .O(new_n677_));
  inv1 g0471(.a(new_n677_), .O(new_n678_));
  nor2 g0472(.a(new_n678_), .b(new_n674_), .O(new_n679_));
  inv1 g0473(.a(new_n679_), .O(o_32_));
  inv1 g0474(.a(i_55_), .O(new_n681_));
  nor2 g0475(.a(new_n504_), .b(new_n681_), .O(new_n682_));
  nor2 g0476(.a(new_n614_), .b(new_n509_), .O(new_n683_));
  nor2 g0477(.a(new_n683_), .b(new_n682_), .O(new_n684_));
  inv1 g0478(.a(new_n684_), .O(o_23_));
  nor2 g0479(.a(new_n634_), .b(new_n478_), .O(new_n686_));
  inv1 g0480(.a(i_52_), .O(new_n687_));
  nor2 g0481(.a(new_n535_), .b(new_n687_), .O(new_n688_));
  nor2 g0482(.a(new_n688_), .b(new_n686_), .O(new_n689_));
  inv1 g0483(.a(new_n689_), .O(o_18_));
  inv1 g0484(.a(i_56_), .O(new_n692_));
  nor2 g0485(.a(new_n504_), .b(new_n692_), .O(new_n693_));
  nor2 g0486(.a(new_n595_), .b(new_n509_), .O(new_n694_));
  nor2 g0487(.a(new_n694_), .b(new_n693_), .O(new_n695_));
  inv1 g0488(.a(new_n695_), .O(o_24_));
  nor2 g0489(.a(new_n634_), .b(new_n492_), .O(new_n697_));
  inv1 g0490(.a(i_51_), .O(new_n698_));
  nor2 g0491(.a(new_n535_), .b(new_n698_), .O(new_n699_));
  nor2 g0492(.a(new_n699_), .b(new_n697_), .O(new_n700_));
  inv1 g0493(.a(new_n700_), .O(o_17_));
  inv1 g0494(.a(i_12_), .O(new_n702_));
  nor2 g0495(.a(i_90_), .b(new_n702_), .O(new_n703_));
  inv1 g0496(.a(i_90_), .O(new_n704_));
  nor2 g0497(.a(new_n704_), .b(i_12_), .O(new_n705_));
  nor2 g0498(.a(new_n705_), .b(new_n703_), .O(new_n706_));
  nor2 g0499(.a(new_n706_), .b(i_82_), .O(new_n707_));
  inv1 g0500(.a(new_n707_), .O(new_n708_));
  nor2 g0501(.a(new_n708_), .b(new_n386_), .O(new_n709_));
  nor2 g0502(.a(new_n706_), .b(i_23_), .O(new_n710_));
  nor2 g0503(.a(new_n376_), .b(i_82_), .O(new_n711_));
  inv1 g0504(.a(new_n711_), .O(new_n712_));
  nor2 g0505(.a(new_n712_), .b(new_n702_), .O(new_n713_));
  nor2 g0506(.a(new_n713_), .b(new_n710_), .O(new_n714_));
  nor2 g0507(.a(i_33_), .b(i_20_), .O(new_n715_));
  inv1 g0508(.a(new_n715_), .O(new_n716_));
  nor2 g0509(.a(new_n716_), .b(new_n714_), .O(new_n717_));
  inv1 g0510(.a(new_n717_), .O(new_n718_));
  nor2 g0511(.a(new_n718_), .b(new_n409_), .O(new_n719_));
  inv1 g0512(.a(i_98_), .O(new_n720_));
  nor2 g0513(.a(new_n428_), .b(new_n720_), .O(new_n721_));
  nor2 g0514(.a(new_n712_), .b(i_12_), .O(new_n722_));
  inv1 g0515(.a(new_n722_), .O(new_n723_));
  nor2 g0516(.a(new_n723_), .b(new_n357_), .O(new_n724_));
  nor2 g0517(.a(new_n724_), .b(new_n377_), .O(new_n725_));
  nor2 g0518(.a(new_n405_), .b(new_n541_), .O(new_n726_));
  inv1 g0519(.a(new_n726_), .O(new_n727_));
  nor2 g0520(.a(new_n727_), .b(new_n725_), .O(new_n728_));
  nor2 g0521(.a(new_n728_), .b(new_n721_), .O(new_n729_));
  inv1 g0522(.a(new_n729_), .O(new_n730_));
  nor2 g0523(.a(new_n730_), .b(new_n719_), .O(new_n731_));
  inv1 g0524(.a(new_n731_), .O(new_n732_));
  nor2 g0525(.a(new_n732_), .b(new_n709_), .O(new_n733_));
  inv1 g0526(.a(new_n733_), .O(o_69_));
  inv1 g0527(.a(i_85_), .O(new_n735_));
  nor2 g0528(.a(new_n451_), .b(new_n735_), .O(new_n736_));
  nor2 g0529(.a(new_n557_), .b(new_n376_), .O(new_n737_));
  inv1 g0530(.a(new_n737_), .O(new_n738_));
  nor2 g0531(.a(new_n738_), .b(new_n407_), .O(new_n739_));
  nor2 g0532(.a(new_n739_), .b(new_n736_), .O(new_n740_));
  inv1 g0533(.a(new_n740_), .O(o_56_));
  inv1 g0534(.a(i_72_), .O(new_n742_));
  nor2 g0535(.a(new_n643_), .b(new_n742_), .O(new_n743_));
  nor2 g0536(.a(new_n646_), .b(new_n275_), .O(new_n744_));
  nor2 g0537(.a(new_n421_), .b(new_n591_), .O(new_n745_));
  inv1 g0538(.a(new_n745_), .O(new_n746_));
  nor2 g0539(.a(new_n746_), .b(new_n482_), .O(new_n747_));
  nor2 g0540(.a(new_n747_), .b(new_n744_), .O(new_n748_));
  inv1 g0541(.a(new_n748_), .O(new_n749_));
  nor2 g0542(.a(new_n749_), .b(new_n743_), .O(new_n750_));
  inv1 g0543(.a(new_n750_), .O(o_43_));
  nor2 g0544(.a(new_n573_), .b(i_22_), .O(new_n753_));
  nor2 g0545(.a(new_n570_), .b(i_84_), .O(new_n754_));
  nor2 g0546(.a(new_n754_), .b(new_n753_), .O(new_n755_));
  nor2 g0547(.a(new_n755_), .b(new_n227_), .O(new_n756_));
  inv1 g0548(.a(new_n756_), .O(o_55_));
  inv1 g0549(.a(i_73_), .O(new_n758_));
  nor2 g0550(.a(new_n643_), .b(new_n758_), .O(new_n759_));
  nor2 g0551(.a(new_n646_), .b(new_n274_), .O(new_n760_));
  nor2 g0552(.a(new_n421_), .b(new_n453_), .O(new_n761_));
  inv1 g0553(.a(new_n761_), .O(new_n762_));
  nor2 g0554(.a(new_n762_), .b(new_n482_), .O(new_n763_));
  nor2 g0555(.a(new_n763_), .b(new_n760_), .O(new_n764_));
  inv1 g0556(.a(new_n764_), .O(new_n765_));
  nor2 g0557(.a(new_n765_), .b(new_n759_), .O(new_n766_));
  inv1 g0558(.a(new_n766_), .O(o_44_));
  inv1 g0559(.a(i_87_), .O(new_n768_));
  nor2 g0560(.a(new_n451_), .b(new_n768_), .O(new_n769_));
  nor2 g0561(.a(new_n454_), .b(new_n572_), .O(new_n770_));
  nor2 g0562(.a(new_n770_), .b(new_n769_), .O(new_n771_));
  inv1 g0563(.a(new_n771_), .O(o_58_));
  inv1 g0564(.a(i_70_), .O(new_n773_));
  nor2 g0565(.a(new_n643_), .b(new_n773_), .O(new_n774_));
  nor2 g0566(.a(new_n646_), .b(new_n271_), .O(new_n775_));
  nor2 g0567(.a(new_n421_), .b(new_n520_), .O(new_n776_));
  inv1 g0568(.a(new_n776_), .O(new_n777_));
  nor2 g0569(.a(new_n777_), .b(new_n482_), .O(new_n778_));
  nor2 g0570(.a(new_n778_), .b(new_n775_), .O(new_n779_));
  inv1 g0571(.a(new_n779_), .O(new_n780_));
  nor2 g0572(.a(new_n780_), .b(new_n774_), .O(new_n781_));
  inv1 g0573(.a(new_n781_), .O(o_41_));
  nor2 g0574(.a(new_n311_), .b(new_n295_), .O(new_n783_));
  inv1 g0575(.a(new_n783_), .O(new_n784_));
  nor2 g0576(.a(new_n784_), .b(new_n267_), .O(new_n785_));
  inv1 g0577(.a(new_n785_), .O(new_n786_));
  nor2 g0578(.a(new_n786_), .b(new_n289_), .O(new_n787_));
  nor2 g0579(.a(new_n333_), .b(new_n311_), .O(new_n788_));
  nor2 g0580(.a(new_n788_), .b(new_n787_), .O(new_n789_));
  nor2 g0581(.a(new_n245_), .b(new_n239_), .O(new_n790_));
  inv1 g0582(.a(new_n790_), .O(new_n791_));
  nor2 g0583(.a(new_n791_), .b(i_108_), .O(new_n792_));
  inv1 g0584(.a(new_n792_), .O(new_n793_));
  nor2 g0585(.a(new_n793_), .b(new_n789_), .O(new_n794_));
  nor2 g0586(.a(new_n323_), .b(new_n256_), .O(new_n795_));
  nor2 g0587(.a(new_n791_), .b(new_n331_), .O(new_n796_));
  nor2 g0588(.a(new_n796_), .b(new_n311_), .O(new_n797_));
  nor2 g0589(.a(new_n797_), .b(new_n795_), .O(new_n798_));
  nor2 g0590(.a(new_n798_), .b(new_n238_), .O(new_n799_));
  nor2 g0591(.a(new_n799_), .b(new_n316_), .O(new_n800_));
  inv1 g0592(.a(new_n800_), .O(new_n801_));
  nor2 g0593(.a(new_n801_), .b(new_n794_), .O(new_n802_));
  inv1 g0594(.a(new_n802_), .O(o_79_));
  inv1 g0595(.a(i_86_), .O(new_n804_));
  nor2 g0596(.a(new_n451_), .b(new_n804_), .O(new_n805_));
  nor2 g0597(.a(new_n520_), .b(new_n376_), .O(new_n806_));
  inv1 g0598(.a(new_n806_), .O(new_n807_));
  nor2 g0599(.a(new_n807_), .b(new_n407_), .O(new_n808_));
  nor2 g0600(.a(new_n808_), .b(new_n805_), .O(new_n809_));
  inv1 g0601(.a(new_n809_), .O(o_57_));
  inv1 g0602(.a(i_71_), .O(new_n811_));
  nor2 g0603(.a(new_n643_), .b(new_n811_), .O(new_n812_));
  nor2 g0604(.a(new_n646_), .b(new_n276_), .O(new_n813_));
  nor2 g0605(.a(new_n421_), .b(new_n572_), .O(new_n814_));
  inv1 g0606(.a(new_n814_), .O(new_n815_));
  nor2 g0607(.a(new_n815_), .b(new_n482_), .O(new_n816_));
  nor2 g0608(.a(new_n816_), .b(new_n813_), .O(new_n817_));
  inv1 g0609(.a(new_n817_), .O(new_n818_));
  nor2 g0610(.a(new_n818_), .b(new_n812_), .O(new_n819_));
  inv1 g0611(.a(new_n819_), .O(o_42_));
  inv1 g0612(.a(i_81_), .O(new_n821_));
  nor2 g0613(.a(new_n570_), .b(new_n821_), .O(new_n822_));
  nor2 g0614(.a(new_n573_), .b(new_n453_), .O(new_n823_));
  nor2 g0615(.a(new_n823_), .b(new_n227_), .O(new_n824_));
  inv1 g0616(.a(new_n824_), .O(new_n825_));
  nor2 g0617(.a(new_n825_), .b(new_n822_), .O(new_n826_));
  inv1 g0618(.a(new_n826_), .O(o_52_));
  inv1 g0619(.a(i_76_), .O(new_n828_));
  nor2 g0620(.a(new_n643_), .b(new_n828_), .O(new_n829_));
  nor2 g0621(.a(new_n646_), .b(new_n279_), .O(new_n830_));
  nor2 g0622(.a(new_n421_), .b(new_n476_), .O(new_n831_));
  inv1 g0623(.a(new_n831_), .O(new_n832_));
  nor2 g0624(.a(new_n832_), .b(new_n482_), .O(new_n833_));
  nor2 g0625(.a(new_n833_), .b(new_n830_), .O(new_n834_));
  inv1 g0626(.a(new_n834_), .O(new_n835_));
  nor2 g0627(.a(new_n835_), .b(new_n829_), .O(new_n836_));
  inv1 g0628(.a(new_n836_), .O(o_47_));
  nor2 g0629(.a(new_n573_), .b(new_n591_), .O(new_n838_));
  inv1 g0630(.a(i_80_), .O(new_n839_));
  nor2 g0631(.a(new_n570_), .b(new_n839_), .O(new_n840_));
  nor2 g0632(.a(new_n840_), .b(new_n227_), .O(new_n841_));
  inv1 g0633(.a(new_n841_), .O(new_n842_));
  nor2 g0634(.a(new_n842_), .b(new_n838_), .O(new_n843_));
  inv1 g0635(.a(new_n843_), .O(o_51_));
  inv1 g0636(.a(i_77_), .O(new_n845_));
  nor2 g0637(.a(new_n570_), .b(new_n845_), .O(new_n846_));
  nor2 g0638(.a(new_n573_), .b(new_n557_), .O(new_n847_));
  nor2 g0639(.a(new_n847_), .b(new_n227_), .O(new_n848_));
  inv1 g0640(.a(new_n848_), .O(new_n849_));
  nor2 g0641(.a(new_n849_), .b(new_n846_), .O(new_n850_));
  inv1 g0642(.a(new_n850_), .O(o_48_));
  inv1 g0643(.a(i_83_), .O(new_n852_));
  nor2 g0644(.a(new_n570_), .b(new_n852_), .O(new_n853_));
  nor2 g0645(.a(new_n573_), .b(new_n430_), .O(new_n854_));
  nor2 g0646(.a(new_n854_), .b(new_n227_), .O(new_n855_));
  inv1 g0647(.a(new_n855_), .O(new_n856_));
  nor2 g0648(.a(new_n856_), .b(new_n853_), .O(new_n857_));
  inv1 g0649(.a(new_n857_), .O(o_54_));
  inv1 g0650(.a(i_74_), .O(new_n859_));
  nor2 g0651(.a(new_n643_), .b(new_n859_), .O(new_n860_));
  nor2 g0652(.a(new_n646_), .b(new_n270_), .O(new_n861_));
  nor2 g0653(.a(new_n421_), .b(new_n541_), .O(new_n862_));
  inv1 g0654(.a(new_n862_), .O(new_n863_));
  nor2 g0655(.a(new_n863_), .b(new_n482_), .O(new_n864_));
  nor2 g0656(.a(new_n864_), .b(new_n861_), .O(new_n865_));
  inv1 g0657(.a(new_n865_), .O(new_n866_));
  nor2 g0658(.a(new_n866_), .b(new_n860_), .O(new_n867_));
  inv1 g0659(.a(new_n867_), .O(o_45_));
  inv1 g0660(.a(i_44_), .O(new_n869_));
  nor2 g0661(.a(new_n369_), .b(new_n361_), .O(new_n870_));
  nor2 g0662(.a(new_n870_), .b(new_n499_), .O(new_n871_));
  nor2 g0663(.a(new_n460_), .b(new_n361_), .O(new_n872_));
  nor2 g0664(.a(new_n359_), .b(new_n373_), .O(new_n873_));
  inv1 g0665(.a(new_n873_), .O(new_n874_));
  nor2 g0666(.a(new_n874_), .b(new_n872_), .O(new_n875_));
  inv1 g0667(.a(new_n875_), .O(new_n876_));
  nor2 g0668(.a(new_n876_), .b(new_n871_), .O(new_n877_));
  nor2 g0669(.a(new_n877_), .b(new_n227_), .O(new_n878_));
  nor2 g0670(.a(new_n368_), .b(new_n515_), .O(new_n879_));
  nor2 g0671(.a(new_n879_), .b(i_26_), .O(new_n880_));
  nor2 g0672(.a(i_24_), .b(i_27_), .O(new_n881_));
  nor2 g0673(.a(new_n881_), .b(new_n227_), .O(new_n882_));
  inv1 g0674(.a(new_n882_), .O(new_n883_));
  nor2 g0675(.a(new_n883_), .b(new_n880_), .O(new_n884_));
  nor2 g0676(.a(new_n884_), .b(new_n878_), .O(new_n885_));
  inv1 g0677(.a(new_n885_), .O(new_n886_));
  inv1 g0678(.a(new_n870_), .O(new_n887_));
  nor2 g0679(.a(new_n887_), .b(new_n227_), .O(new_n888_));
  nor2 g0680(.a(new_n888_), .b(new_n886_), .O(new_n889_));
  nor2 g0681(.a(new_n889_), .b(new_n869_), .O(new_n890_));
  inv1 g0682(.a(new_n470_), .O(new_n891_));
  nor2 g0683(.a(new_n891_), .b(new_n458_), .O(new_n892_));
  nor2 g0684(.a(new_n530_), .b(new_n469_), .O(new_n893_));
  inv1 g0685(.a(new_n893_), .O(new_n894_));
  nor2 g0686(.a(new_n894_), .b(new_n687_), .O(new_n895_));
  nor2 g0687(.a(new_n895_), .b(new_n892_), .O(new_n896_));
  inv1 g0688(.a(new_n896_), .O(new_n897_));
  inv1 g0689(.a(new_n642_), .O(new_n898_));
  nor2 g0690(.a(new_n898_), .b(new_n828_), .O(new_n899_));
  inv1 g0691(.a(i_84_), .O(new_n900_));
  nor2 g0692(.a(new_n375_), .b(new_n363_), .O(new_n901_));
  inv1 g0693(.a(new_n901_), .O(new_n902_));
  nor2 g0694(.a(new_n902_), .b(new_n569_), .O(new_n903_));
  inv1 g0695(.a(new_n903_), .O(new_n904_));
  nor2 g0696(.a(new_n904_), .b(new_n900_), .O(new_n905_));
  nor2 g0697(.a(new_n905_), .b(new_n899_), .O(new_n906_));
  inv1 g0698(.a(new_n906_), .O(new_n907_));
  inv1 g0699(.a(i_100_), .O(new_n908_));
  nor2 g0700(.a(new_n902_), .b(new_n423_), .O(new_n909_));
  inv1 g0701(.a(new_n909_), .O(new_n910_));
  nor2 g0702(.a(new_n910_), .b(new_n908_), .O(new_n911_));
  inv1 g0703(.a(i_92_), .O(new_n912_));
  nor2 g0704(.a(new_n567_), .b(new_n376_), .O(new_n913_));
  inv1 g0705(.a(new_n913_), .O(new_n914_));
  nor2 g0706(.a(new_n914_), .b(new_n902_), .O(new_n915_));
  inv1 g0707(.a(new_n915_), .O(new_n916_));
  nor2 g0708(.a(new_n916_), .b(new_n912_), .O(new_n917_));
  nor2 g0709(.a(new_n917_), .b(new_n911_), .O(new_n918_));
  inv1 g0710(.a(new_n918_), .O(new_n919_));
  nor2 g0711(.a(new_n919_), .b(new_n907_), .O(new_n920_));
  inv1 g0712(.a(new_n920_), .O(new_n921_));
  nor2 g0713(.a(new_n921_), .b(new_n897_), .O(new_n922_));
  inv1 g0714(.a(new_n922_), .O(new_n923_));
  nor2 g0715(.a(new_n923_), .b(new_n890_), .O(new_n924_));
  inv1 g0716(.a(new_n924_), .O(o_10_));
  inv1 g0717(.a(i_82_), .O(new_n926_));
  nor2 g0718(.a(new_n570_), .b(new_n926_), .O(new_n927_));
  nor2 g0719(.a(new_n573_), .b(new_n541_), .O(new_n928_));
  nor2 g0720(.a(new_n928_), .b(new_n227_), .O(new_n929_));
  inv1 g0721(.a(new_n929_), .O(new_n930_));
  nor2 g0722(.a(new_n930_), .b(new_n927_), .O(new_n931_));
  inv1 g0723(.a(new_n931_), .O(o_53_));
  inv1 g0724(.a(i_75_), .O(new_n933_));
  nor2 g0725(.a(new_n643_), .b(new_n933_), .O(new_n934_));
  nor2 g0726(.a(new_n646_), .b(new_n280_), .O(new_n935_));
  inv1 g0727(.a(new_n431_), .O(new_n936_));
  nor2 g0728(.a(new_n482_), .b(new_n936_), .O(new_n937_));
  nor2 g0729(.a(new_n937_), .b(new_n935_), .O(new_n938_));
  inv1 g0730(.a(new_n938_), .O(new_n939_));
  nor2 g0731(.a(new_n939_), .b(new_n934_), .O(new_n940_));
  inv1 g0732(.a(new_n940_), .O(o_46_));
  nor2 g0733(.a(new_n274_), .b(new_n270_), .O(new_n942_));
  inv1 g0734(.a(new_n942_), .O(new_n943_));
  nor2 g0735(.a(new_n305_), .b(new_n278_), .O(new_n944_));
  inv1 g0736(.a(new_n944_), .O(new_n945_));
  nor2 g0737(.a(new_n945_), .b(new_n786_), .O(new_n946_));
  nor2 g0738(.a(new_n946_), .b(new_n788_), .O(new_n947_));
  nor2 g0739(.a(new_n947_), .b(new_n943_), .O(new_n948_));
  inv1 g0740(.a(new_n948_), .O(new_n949_));
  nor2 g0741(.a(new_n280_), .b(i_116_), .O(new_n950_));
  inv1 g0742(.a(new_n950_), .O(new_n951_));
  nor2 g0743(.a(new_n951_), .b(new_n949_), .O(new_n952_));
  nor2 g0744(.a(new_n247_), .b(new_n248_), .O(new_n953_));
  nor2 g0745(.a(new_n953_), .b(new_n321_), .O(new_n954_));
  nor2 g0746(.a(i_33_), .b(new_n280_), .O(new_n955_));
  inv1 g0747(.a(new_n955_), .O(new_n956_));
  nor2 g0748(.a(new_n956_), .b(new_n943_), .O(new_n957_));
  inv1 g0749(.a(new_n957_), .O(new_n958_));
  nor2 g0750(.a(new_n958_), .b(new_n954_), .O(new_n959_));
  nor2 g0751(.a(new_n959_), .b(new_n311_), .O(new_n960_));
  nor2 g0752(.a(new_n311_), .b(new_n234_), .O(new_n961_));
  nor2 g0753(.a(new_n303_), .b(new_n278_), .O(new_n962_));
  inv1 g0754(.a(new_n962_), .O(new_n963_));
  nor2 g0755(.a(new_n963_), .b(new_n255_), .O(new_n964_));
  nor2 g0756(.a(new_n964_), .b(new_n323_), .O(new_n965_));
  nor2 g0757(.a(new_n965_), .b(new_n961_), .O(new_n966_));
  inv1 g0758(.a(new_n966_), .O(new_n967_));
  nor2 g0759(.a(new_n967_), .b(new_n960_), .O(new_n968_));
  nor2 g0760(.a(new_n968_), .b(new_n279_), .O(new_n969_));
  nor2 g0761(.a(new_n969_), .b(new_n316_), .O(new_n970_));
  inv1 g0762(.a(new_n970_), .O(new_n971_));
  nor2 g0763(.a(new_n971_), .b(new_n952_), .O(new_n972_));
  inv1 g0764(.a(new_n972_), .O(o_87_));
  nor2 g0765(.a(new_n786_), .b(i_102_), .O(new_n974_));
  nor2 g0766(.a(new_n785_), .b(new_n311_), .O(new_n975_));
  nor2 g0767(.a(new_n975_), .b(new_n974_), .O(new_n976_));
  nor2 g0768(.a(new_n976_), .b(new_n251_), .O(new_n977_));
  nor2 g0769(.a(i_103_), .b(new_n250_), .O(new_n978_));
  inv1 g0770(.a(new_n978_), .O(new_n979_));
  nor2 g0771(.a(new_n979_), .b(new_n786_), .O(new_n980_));
  nor2 g0772(.a(new_n980_), .b(new_n316_), .O(new_n981_));
  inv1 g0773(.a(new_n981_), .O(new_n982_));
  nor2 g0774(.a(new_n982_), .b(new_n977_), .O(new_n983_));
  inv1 g0775(.a(new_n983_), .O(o_74_));
  nor2 g0776(.a(new_n451_), .b(new_n704_), .O(new_n985_));
  nor2 g0777(.a(new_n454_), .b(new_n541_), .O(new_n986_));
  nor2 g0778(.a(new_n986_), .b(new_n985_), .O(new_n987_));
  inv1 g0779(.a(new_n987_), .O(o_61_));
  inv1 g0780(.a(i_43_), .O(new_n989_));
  nor2 g0781(.a(new_n889_), .b(new_n989_), .O(new_n990_));
  nor2 g0782(.a(new_n891_), .b(new_n488_), .O(new_n991_));
  nor2 g0783(.a(new_n894_), .b(new_n698_), .O(new_n992_));
  nor2 g0784(.a(new_n992_), .b(new_n991_), .O(new_n993_));
  inv1 g0785(.a(new_n993_), .O(new_n994_));
  nor2 g0786(.a(new_n898_), .b(new_n933_), .O(new_n995_));
  nor2 g0787(.a(new_n904_), .b(new_n852_), .O(new_n996_));
  nor2 g0788(.a(new_n996_), .b(new_n995_), .O(new_n997_));
  inv1 g0789(.a(new_n997_), .O(new_n998_));
  nor2 g0790(.a(new_n910_), .b(new_n420_), .O(new_n999_));
  nor2 g0791(.a(new_n916_), .b(new_n388_), .O(new_n1000_));
  nor2 g0792(.a(new_n1000_), .b(new_n999_), .O(new_n1001_));
  inv1 g0793(.a(new_n1001_), .O(new_n1002_));
  nor2 g0794(.a(new_n1002_), .b(new_n998_), .O(new_n1003_));
  inv1 g0795(.a(new_n1003_), .O(new_n1004_));
  nor2 g0796(.a(new_n1004_), .b(new_n994_), .O(new_n1005_));
  inv1 g0797(.a(new_n1005_), .O(new_n1006_));
  nor2 g0798(.a(new_n1006_), .b(new_n990_), .O(new_n1007_));
  inv1 g0799(.a(new_n1007_), .O(o_9_));
  inv1 g0800(.a(new_n975_), .O(new_n1009_));
  nor2 g0801(.a(new_n1009_), .b(new_n250_), .O(new_n1010_));
  nor2 g0802(.a(new_n974_), .b(new_n316_), .O(new_n1011_));
  inv1 g0803(.a(new_n1011_), .O(new_n1012_));
  nor2 g0804(.a(new_n1012_), .b(new_n1010_), .O(new_n1013_));
  inv1 g0805(.a(new_n1013_), .O(o_73_));
  nor2 g0806(.a(new_n451_), .b(new_n388_), .O(new_n1015_));
  nor2 g0807(.a(new_n433_), .b(new_n407_), .O(new_n1016_));
  nor2 g0808(.a(new_n1016_), .b(new_n1015_), .O(new_n1017_));
  inv1 g0809(.a(new_n1017_), .O(o_62_));
  nor2 g0810(.a(new_n943_), .b(new_n331_), .O(new_n1019_));
  nor2 g0811(.a(new_n1019_), .b(new_n311_), .O(new_n1020_));
  nor2 g0812(.a(new_n965_), .b(new_n324_), .O(new_n1021_));
  inv1 g0813(.a(new_n1021_), .O(new_n1022_));
  nor2 g0814(.a(new_n1022_), .b(new_n1020_), .O(new_n1023_));
  nor2 g0815(.a(new_n1023_), .b(new_n270_), .O(new_n1024_));
  nor2 g0816(.a(new_n274_), .b(i_114_), .O(new_n1025_));
  inv1 g0817(.a(new_n1025_), .O(new_n1026_));
  nor2 g0818(.a(new_n1026_), .b(new_n947_), .O(new_n1027_));
  nor2 g0819(.a(new_n1027_), .b(new_n316_), .O(new_n1028_));
  inv1 g0820(.a(new_n1028_), .O(new_n1029_));
  nor2 g0821(.a(new_n1029_), .b(new_n1024_), .O(new_n1030_));
  inv1 g0822(.a(new_n1030_), .O(o_85_));
  nor2 g0823(.a(new_n305_), .b(new_n336_), .O(new_n1032_));
  nor2 g0824(.a(new_n1032_), .b(new_n269_), .O(new_n1033_));
  nor2 g0825(.a(i_101_), .b(new_n227_), .O(new_n1034_));
  inv1 g0826(.a(new_n1034_), .O(new_n1035_));
  nor2 g0827(.a(new_n1035_), .b(new_n267_), .O(new_n1036_));
  nor2 g0828(.a(new_n1036_), .b(new_n1033_), .O(new_n1037_));
  nor2 g0829(.a(new_n1037_), .b(new_n293_), .O(new_n1038_));
  inv1 g0830(.a(new_n325_), .O(new_n1039_));
  nor2 g0831(.a(new_n1039_), .b(new_n249_), .O(new_n1040_));
  nor2 g0832(.a(new_n1040_), .b(new_n316_), .O(new_n1041_));
  inv1 g0833(.a(new_n1041_), .O(new_n1042_));
  nor2 g0834(.a(new_n1042_), .b(new_n1038_), .O(new_n1043_));
  inv1 g0835(.a(new_n1043_), .O(o_72_));
  nor2 g0836(.a(new_n451_), .b(new_n912_), .O(new_n1045_));
  nor2 g0837(.a(new_n454_), .b(new_n476_), .O(new_n1046_));
  nor2 g0838(.a(new_n1046_), .b(new_n1045_), .O(new_n1047_));
  inv1 g0839(.a(new_n1047_), .O(o_63_));
  inv1 g0840(.a(i_78_), .O(new_n1049_));
  nor2 g0841(.a(new_n570_), .b(new_n1049_), .O(new_n1050_));
  nor2 g0842(.a(new_n573_), .b(new_n520_), .O(new_n1051_));
  nor2 g0843(.a(new_n1051_), .b(new_n227_), .O(new_n1052_));
  inv1 g0844(.a(new_n1052_), .O(new_n1053_));
  nor2 g0845(.a(new_n1053_), .b(new_n1050_), .O(new_n1054_));
  inv1 g0846(.a(new_n1054_), .O(o_49_));
  inv1 g0847(.a(new_n888_), .O(new_n1056_));
  nor2 g0848(.a(new_n1056_), .b(new_n876_), .O(new_n1057_));
  inv1 g0849(.a(new_n1057_), .O(new_n1058_));
  nor2 g0850(.a(new_n1058_), .b(new_n498_), .O(new_n1059_));
  nor2 g0851(.a(new_n916_), .b(new_n448_), .O(new_n1060_));
  inv1 g0852(.a(i_41_), .O(new_n1061_));
  inv1 g0853(.a(new_n884_), .O(new_n1062_));
  nor2 g0854(.a(new_n1062_), .b(new_n1061_), .O(new_n1063_));
  nor2 g0855(.a(new_n1063_), .b(new_n1060_), .O(new_n1064_));
  inv1 g0856(.a(new_n1064_), .O(new_n1065_));
  nor2 g0857(.a(new_n904_), .b(new_n821_), .O(new_n1066_));
  nor2 g0858(.a(new_n894_), .b(new_n668_), .O(new_n1067_));
  nor2 g0859(.a(new_n1067_), .b(new_n1066_), .O(new_n1068_));
  inv1 g0860(.a(new_n1068_), .O(new_n1069_));
  nor2 g0861(.a(new_n1069_), .b(new_n1065_), .O(new_n1070_));
  inv1 g0862(.a(new_n1070_), .O(new_n1071_));
  nor2 g0863(.a(new_n1071_), .b(new_n1059_), .O(new_n1072_));
  inv1 g0864(.a(new_n1072_), .O(new_n1073_));
  inv1 g0865(.a(new_n878_), .O(new_n1074_));
  nor2 g0866(.a(new_n1074_), .b(new_n1061_), .O(new_n1075_));
  nor2 g0867(.a(new_n898_), .b(new_n758_), .O(new_n1076_));
  nor2 g0868(.a(new_n891_), .b(new_n579_), .O(new_n1077_));
  inv1 g0869(.a(i_97_), .O(new_n1078_));
  nor2 g0870(.a(new_n910_), .b(new_n1078_), .O(new_n1079_));
  nor2 g0871(.a(new_n1079_), .b(new_n1077_), .O(new_n1080_));
  inv1 g0872(.a(new_n1080_), .O(new_n1081_));
  nor2 g0873(.a(new_n1081_), .b(new_n1076_), .O(new_n1082_));
  inv1 g0874(.a(new_n1082_), .O(new_n1083_));
  nor2 g0875(.a(new_n1083_), .b(new_n1075_), .O(new_n1084_));
  inv1 g0876(.a(new_n1084_), .O(new_n1085_));
  nor2 g0877(.a(new_n1085_), .b(new_n1073_), .O(new_n1086_));
  inv1 g0878(.a(new_n1086_), .O(o_7_));
  nor2 g0879(.a(new_n949_), .b(i_115_), .O(new_n1088_));
  nor2 g0880(.a(new_n1023_), .b(new_n280_), .O(new_n1089_));
  nor2 g0881(.a(new_n1089_), .b(new_n316_), .O(new_n1090_));
  inv1 g0882(.a(new_n1090_), .O(new_n1091_));
  nor2 g0883(.a(new_n1091_), .b(new_n1088_), .O(new_n1092_));
  inv1 g0884(.a(new_n1092_), .O(o_86_));
  inv1 g0885(.a(new_n364_), .O(new_n1094_));
  nor2 g0886(.a(new_n379_), .b(new_n368_), .O(new_n1095_));
  inv1 g0887(.a(new_n1095_), .O(new_n1096_));
  nor2 g0888(.a(new_n1096_), .b(new_n1094_), .O(new_n1097_));
  nor2 g0889(.a(new_n1097_), .b(i_84_), .O(new_n1098_));
  nor2 g0890(.a(new_n1098_), .b(new_n753_), .O(new_n1099_));
  inv1 g0891(.a(i_14_), .O(new_n1100_));
  nor2 g0892(.a(new_n227_), .b(new_n1100_), .O(new_n1101_));
  inv1 g0893(.a(new_n1101_), .O(new_n1102_));
  nor2 g0894(.a(new_n1102_), .b(new_n357_), .O(new_n1103_));
  inv1 g0895(.a(new_n1103_), .O(new_n1104_));
  nor2 g0896(.a(new_n1104_), .b(new_n1099_), .O(new_n1105_));
  nor2 g0897(.a(new_n428_), .b(new_n908_), .O(new_n1106_));
  nor2 g0898(.a(new_n832_), .b(new_n405_), .O(new_n1107_));
  nor2 g0899(.a(new_n1107_), .b(new_n1106_), .O(new_n1108_));
  inv1 g0900(.a(new_n1108_), .O(new_n1109_));
  nor2 g0901(.a(new_n1109_), .b(new_n1105_), .O(new_n1110_));
  inv1 g0902(.a(new_n1110_), .O(o_71_));
  nor2 g0903(.a(i_7_), .b(i_85_), .O(new_n1112_));
  inv1 g0904(.a(i_7_), .O(new_n1113_));
  nor2 g0905(.a(new_n1113_), .b(new_n735_), .O(new_n1114_));
  nor2 g0906(.a(new_n1114_), .b(new_n1112_), .O(new_n1115_));
  inv1 g0907(.a(new_n1115_), .O(new_n1116_));
  nor2 g0908(.a(new_n1116_), .b(i_77_), .O(new_n1117_));
  inv1 g0909(.a(new_n1117_), .O(new_n1118_));
  nor2 g0910(.a(new_n1118_), .b(new_n386_), .O(new_n1119_));
  nor2 g0911(.a(new_n1116_), .b(i_23_), .O(new_n1120_));
  nor2 g0912(.a(new_n376_), .b(i_77_), .O(new_n1121_));
  inv1 g0913(.a(new_n1121_), .O(new_n1122_));
  nor2 g0914(.a(new_n1122_), .b(new_n1113_), .O(new_n1123_));
  nor2 g0915(.a(new_n1123_), .b(new_n1120_), .O(new_n1124_));
  nor2 g0916(.a(i_33_), .b(i_15_), .O(new_n1125_));
  inv1 g0917(.a(new_n1125_), .O(new_n1126_));
  nor2 g0918(.a(new_n1126_), .b(new_n1124_), .O(new_n1127_));
  inv1 g0919(.a(new_n1127_), .O(new_n1128_));
  nor2 g0920(.a(new_n1128_), .b(new_n409_), .O(new_n1129_));
  nor2 g0921(.a(new_n557_), .b(i_7_), .O(new_n1130_));
  inv1 g0922(.a(new_n1130_), .O(new_n1131_));
  nor2 g0923(.a(new_n1131_), .b(new_n1122_), .O(new_n1132_));
  inv1 g0924(.a(new_n1132_), .O(new_n1133_));
  nor2 g0925(.a(new_n1133_), .b(new_n357_), .O(new_n1134_));
  nor2 g0926(.a(new_n1134_), .b(new_n648_), .O(new_n1135_));
  nor2 g0927(.a(new_n1135_), .b(new_n405_), .O(new_n1136_));
  inv1 g0928(.a(i_93_), .O(new_n1137_));
  nor2 g0929(.a(new_n428_), .b(new_n1137_), .O(new_n1138_));
  nor2 g0930(.a(new_n1138_), .b(new_n1136_), .O(new_n1139_));
  inv1 g0931(.a(new_n1139_), .O(new_n1140_));
  nor2 g0932(.a(new_n1140_), .b(new_n1129_), .O(new_n1141_));
  inv1 g0933(.a(new_n1141_), .O(new_n1142_));
  nor2 g0934(.a(new_n1142_), .b(new_n1119_), .O(new_n1143_));
  inv1 g0935(.a(new_n1143_), .O(o_64_));
  inv1 g0936(.a(i_42_), .O(new_n1145_));
  nor2 g0937(.a(new_n885_), .b(new_n1145_), .O(new_n1146_));
  nor2 g0938(.a(new_n891_), .b(new_n539_), .O(new_n1147_));
  nor2 g0939(.a(new_n898_), .b(new_n859_), .O(new_n1148_));
  nor2 g0940(.a(new_n1148_), .b(new_n1147_), .O(new_n1149_));
  inv1 g0941(.a(new_n1149_), .O(new_n1150_));
  nor2 g0942(.a(new_n916_), .b(new_n704_), .O(new_n1151_));
  nor2 g0943(.a(new_n904_), .b(new_n926_), .O(new_n1152_));
  nor2 g0944(.a(new_n1152_), .b(new_n1151_), .O(new_n1153_));
  inv1 g0945(.a(new_n1153_), .O(new_n1154_));
  nor2 g0946(.a(new_n1154_), .b(new_n1150_), .O(new_n1155_));
  inv1 g0947(.a(new_n1155_), .O(new_n1156_));
  nor2 g0948(.a(new_n1058_), .b(new_n551_), .O(new_n1157_));
  nor2 g0949(.a(new_n910_), .b(new_n720_), .O(new_n1158_));
  nor2 g0950(.a(new_n894_), .b(new_n631_), .O(new_n1159_));
  nor2 g0951(.a(new_n1159_), .b(new_n1158_), .O(new_n1160_));
  inv1 g0952(.a(new_n1160_), .O(new_n1161_));
  nor2 g0953(.a(new_n1161_), .b(new_n1157_), .O(new_n1162_));
  inv1 g0954(.a(new_n1162_), .O(new_n1163_));
  nor2 g0955(.a(new_n1163_), .b(new_n1156_), .O(new_n1164_));
  inv1 g0956(.a(new_n1164_), .O(new_n1165_));
  nor2 g0957(.a(new_n1165_), .b(new_n1146_), .O(new_n1166_));
  inv1 g0958(.a(new_n1166_), .O(o_8_));
  inv1 g0959(.a(new_n787_), .O(new_n1168_));
  nor2 g0960(.a(new_n1168_), .b(new_n247_), .O(new_n1169_));
  nor2 g0961(.a(new_n1169_), .b(new_n788_), .O(new_n1170_));
  nor2 g0962(.a(new_n1170_), .b(new_n303_), .O(new_n1171_));
  inv1 g0963(.a(new_n1171_), .O(new_n1172_));
  nor2 g0964(.a(new_n276_), .b(i_112_), .O(new_n1173_));
  inv1 g0965(.a(new_n1173_), .O(new_n1174_));
  nor2 g0966(.a(new_n1174_), .b(new_n1172_), .O(new_n1175_));
  nor2 g0967(.a(new_n254_), .b(new_n321_), .O(new_n1176_));
  nor2 g0968(.a(new_n276_), .b(new_n220_), .O(new_n1177_));
  inv1 g0969(.a(new_n1177_), .O(new_n1178_));
  nor2 g0970(.a(new_n1178_), .b(new_n303_), .O(new_n1179_));
  inv1 g0971(.a(new_n1179_), .O(new_n1180_));
  nor2 g0972(.a(new_n1180_), .b(new_n357_), .O(new_n1181_));
  inv1 g0973(.a(new_n1181_), .O(new_n1182_));
  nor2 g0974(.a(new_n1182_), .b(new_n1176_), .O(new_n1183_));
  inv1 g0975(.a(new_n1183_), .O(new_n1184_));
  nor2 g0976(.a(new_n1184_), .b(new_n954_), .O(new_n1185_));
  nor2 g0977(.a(new_n311_), .b(new_n275_), .O(new_n1186_));
  inv1 g0978(.a(new_n1186_), .O(new_n1187_));
  nor2 g0979(.a(new_n1187_), .b(new_n1185_), .O(new_n1188_));
  nor2 g0980(.a(new_n1188_), .b(new_n316_), .O(new_n1189_));
  inv1 g0981(.a(new_n1189_), .O(new_n1190_));
  nor2 g0982(.a(new_n1190_), .b(new_n1175_), .O(new_n1191_));
  inv1 g0983(.a(new_n1191_), .O(o_83_));
  nor2 g0984(.a(new_n245_), .b(i_107_), .O(new_n1193_));
  inv1 g0985(.a(new_n1193_), .O(new_n1194_));
  nor2 g0986(.a(new_n1194_), .b(new_n789_), .O(new_n1195_));
  nor2 g0987(.a(new_n798_), .b(new_n239_), .O(new_n1196_));
  nor2 g0988(.a(new_n1196_), .b(new_n316_), .O(new_n1197_));
  inv1 g0989(.a(new_n1197_), .O(new_n1198_));
  nor2 g0990(.a(new_n1198_), .b(new_n1195_), .O(new_n1199_));
  inv1 g0991(.a(new_n1199_), .O(o_78_));
  nor2 g0992(.a(i_8_), .b(i_86_), .O(new_n1201_));
  inv1 g0993(.a(i_8_), .O(new_n1202_));
  nor2 g0994(.a(new_n1202_), .b(new_n804_), .O(new_n1203_));
  nor2 g0995(.a(new_n1203_), .b(new_n1201_), .O(new_n1204_));
  inv1 g0996(.a(new_n1204_), .O(new_n1205_));
  nor2 g0997(.a(new_n1205_), .b(i_78_), .O(new_n1206_));
  inv1 g0998(.a(new_n1206_), .O(new_n1207_));
  nor2 g0999(.a(new_n1207_), .b(new_n386_), .O(new_n1208_));
  nor2 g1000(.a(new_n1205_), .b(i_23_), .O(new_n1209_));
  nor2 g1001(.a(new_n376_), .b(i_78_), .O(new_n1210_));
  inv1 g1002(.a(new_n1210_), .O(new_n1211_));
  nor2 g1003(.a(new_n1211_), .b(new_n1202_), .O(new_n1212_));
  nor2 g1004(.a(new_n1212_), .b(new_n1209_), .O(new_n1213_));
  nor2 g1005(.a(i_33_), .b(i_16_), .O(new_n1214_));
  inv1 g1006(.a(new_n1214_), .O(new_n1215_));
  nor2 g1007(.a(new_n1215_), .b(new_n1213_), .O(new_n1216_));
  inv1 g1008(.a(new_n1216_), .O(new_n1217_));
  nor2 g1009(.a(new_n1217_), .b(new_n409_), .O(new_n1218_));
  nor2 g1010(.a(new_n520_), .b(i_8_), .O(new_n1219_));
  inv1 g1011(.a(new_n1219_), .O(new_n1220_));
  nor2 g1012(.a(new_n1220_), .b(new_n1211_), .O(new_n1221_));
  inv1 g1013(.a(new_n1221_), .O(new_n1222_));
  nor2 g1014(.a(new_n1222_), .b(new_n357_), .O(new_n1223_));
  nor2 g1015(.a(new_n1223_), .b(new_n776_), .O(new_n1224_));
  nor2 g1016(.a(new_n1224_), .b(new_n405_), .O(new_n1225_));
  inv1 g1017(.a(i_94_), .O(new_n1226_));
  nor2 g1018(.a(new_n428_), .b(new_n1226_), .O(new_n1227_));
  nor2 g1019(.a(new_n1227_), .b(new_n1225_), .O(new_n1228_));
  inv1 g1020(.a(new_n1228_), .O(new_n1229_));
  nor2 g1021(.a(new_n1229_), .b(new_n1218_), .O(new_n1230_));
  inv1 g1022(.a(new_n1230_), .O(new_n1231_));
  nor2 g1023(.a(new_n1231_), .b(new_n1208_), .O(new_n1232_));
  inv1 g1024(.a(new_n1232_), .O(o_65_));
  inv1 g1025(.a(i_39_), .O(new_n1234_));
  nor2 g1026(.a(new_n885_), .b(new_n1234_), .O(new_n1235_));
  nor2 g1027(.a(new_n891_), .b(new_n618_), .O(new_n1236_));
  nor2 g1028(.a(new_n898_), .b(new_n811_), .O(new_n1237_));
  nor2 g1029(.a(new_n1237_), .b(new_n1236_), .O(new_n1238_));
  inv1 g1030(.a(new_n1238_), .O(new_n1239_));
  nor2 g1031(.a(new_n916_), .b(new_n768_), .O(new_n1240_));
  nor2 g1032(.a(new_n904_), .b(new_n565_), .O(new_n1241_));
  nor2 g1033(.a(new_n1241_), .b(new_n1240_), .O(new_n1242_));
  inv1 g1034(.a(new_n1242_), .O(new_n1243_));
  nor2 g1035(.a(new_n1243_), .b(new_n1239_), .O(new_n1244_));
  inv1 g1036(.a(new_n1244_), .O(new_n1245_));
  nor2 g1037(.a(new_n1058_), .b(new_n681_), .O(new_n1246_));
  inv1 g1038(.a(i_95_), .O(new_n1247_));
  nor2 g1039(.a(new_n910_), .b(new_n1247_), .O(new_n1248_));
  nor2 g1040(.a(new_n894_), .b(new_n609_), .O(new_n1249_));
  nor2 g1041(.a(new_n1249_), .b(new_n1248_), .O(new_n1250_));
  inv1 g1042(.a(new_n1250_), .O(new_n1251_));
  nor2 g1043(.a(new_n1251_), .b(new_n1246_), .O(new_n1252_));
  inv1 g1044(.a(new_n1252_), .O(new_n1253_));
  nor2 g1045(.a(new_n1253_), .b(new_n1245_), .O(new_n1254_));
  inv1 g1046(.a(new_n1254_), .O(new_n1255_));
  nor2 g1047(.a(new_n1255_), .b(new_n1235_), .O(new_n1256_));
  inv1 g1048(.a(new_n1256_), .O(o_5_));
  nor2 g1049(.a(new_n946_), .b(new_n339_), .O(new_n1258_));
  nor2 g1050(.a(new_n1258_), .b(i_113_), .O(new_n1259_));
  nor2 g1051(.a(new_n964_), .b(new_n321_), .O(new_n1260_));
  nor2 g1052(.a(new_n1260_), .b(new_n329_), .O(new_n1261_));
  nor2 g1053(.a(new_n1261_), .b(new_n313_), .O(new_n1262_));
  nor2 g1054(.a(new_n1262_), .b(new_n316_), .O(new_n1263_));
  inv1 g1055(.a(new_n1263_), .O(new_n1264_));
  nor2 g1056(.a(new_n954_), .b(new_n226_), .O(new_n1265_));
  nor2 g1057(.a(new_n1265_), .b(new_n313_), .O(new_n1266_));
  nor2 g1058(.a(new_n335_), .b(new_n308_), .O(new_n1267_));
  nor2 g1059(.a(new_n335_), .b(new_n272_), .O(new_n1268_));
  nor2 g1060(.a(new_n1268_), .b(new_n1267_), .O(new_n1269_));
  inv1 g1061(.a(new_n1269_), .O(new_n1270_));
  nor2 g1062(.a(new_n1270_), .b(new_n1266_), .O(new_n1271_));
  inv1 g1063(.a(new_n1271_), .O(new_n1272_));
  nor2 g1064(.a(new_n1272_), .b(new_n1264_), .O(new_n1273_));
  inv1 g1065(.a(new_n1273_), .O(new_n1274_));
  nor2 g1066(.a(new_n1274_), .b(new_n1259_), .O(new_n1275_));
  inv1 g1067(.a(new_n1275_), .O(o_84_));
  nor2 g1068(.a(new_n243_), .b(i_106_), .O(new_n1277_));
  inv1 g1069(.a(new_n1277_), .O(new_n1278_));
  nor2 g1070(.a(new_n1278_), .b(new_n789_), .O(new_n1279_));
  nor2 g1071(.a(new_n795_), .b(new_n243_), .O(new_n1280_));
  inv1 g1072(.a(new_n1280_), .O(new_n1281_));
  nor2 g1073(.a(new_n1281_), .b(new_n325_), .O(new_n1282_));
  nor2 g1074(.a(new_n311_), .b(new_n242_), .O(new_n1283_));
  inv1 g1075(.a(new_n1283_), .O(new_n1284_));
  nor2 g1076(.a(new_n1284_), .b(new_n1282_), .O(new_n1285_));
  nor2 g1077(.a(new_n1285_), .b(new_n316_), .O(new_n1286_));
  inv1 g1078(.a(new_n1286_), .O(new_n1287_));
  nor2 g1079(.a(new_n1287_), .b(new_n1279_), .O(new_n1288_));
  inv1 g1080(.a(new_n1288_), .O(o_77_));
  nor2 g1081(.a(new_n428_), .b(new_n1247_), .O(new_n1290_));
  inv1 g1082(.a(i_9_), .O(new_n1291_));
  nor2 g1083(.a(i_79_), .b(new_n1291_), .O(new_n1292_));
  inv1 g1084(.a(new_n1292_), .O(new_n1293_));
  nor2 g1085(.a(new_n1293_), .b(new_n227_), .O(new_n1294_));
  inv1 g1086(.a(new_n1294_), .O(new_n1295_));
  nor2 g1087(.a(new_n1295_), .b(new_n357_), .O(new_n1296_));
  inv1 g1088(.a(new_n1296_), .O(new_n1297_));
  nor2 g1089(.a(new_n1297_), .b(new_n1097_), .O(new_n1298_));
  nor2 g1090(.a(new_n815_), .b(new_n405_), .O(new_n1299_));
  nor2 g1091(.a(i_28_), .b(i_27_), .O(new_n1300_));
  inv1 g1092(.a(new_n1300_), .O(new_n1301_));
  nor2 g1093(.a(new_n1301_), .b(new_n357_), .O(new_n1302_));
  inv1 g1094(.a(new_n1302_), .O(new_n1303_));
  nor2 g1095(.a(new_n352_), .b(i_26_), .O(new_n1304_));
  inv1 g1096(.a(new_n1304_), .O(new_n1305_));
  nor2 g1097(.a(i_23_), .b(new_n1291_), .O(new_n1306_));
  inv1 g1098(.a(new_n1306_), .O(new_n1307_));
  nor2 g1099(.a(new_n1307_), .b(i_17_), .O(new_n1308_));
  inv1 g1100(.a(new_n1308_), .O(new_n1309_));
  nor2 g1101(.a(new_n1309_), .b(new_n567_), .O(new_n1310_));
  inv1 g1102(.a(new_n1310_), .O(new_n1311_));
  nor2 g1103(.a(new_n1311_), .b(new_n1305_), .O(new_n1312_));
  inv1 g1104(.a(new_n1312_), .O(new_n1313_));
  nor2 g1105(.a(new_n1313_), .b(new_n1303_), .O(new_n1314_));
  nor2 g1106(.a(new_n1314_), .b(new_n1299_), .O(new_n1315_));
  inv1 g1107(.a(new_n1315_), .O(new_n1316_));
  nor2 g1108(.a(new_n1316_), .b(new_n1298_), .O(new_n1317_));
  inv1 g1109(.a(new_n1317_), .O(new_n1318_));
  nor2 g1110(.a(new_n1318_), .b(new_n1290_), .O(new_n1319_));
  inv1 g1111(.a(new_n1319_), .O(o_66_));
  inv1 g1112(.a(i_88_), .O(new_n1321_));
  nor2 g1113(.a(new_n451_), .b(new_n1321_), .O(new_n1322_));
  nor2 g1114(.a(new_n454_), .b(new_n591_), .O(new_n1323_));
  nor2 g1115(.a(new_n1323_), .b(new_n1322_), .O(new_n1324_));
  inv1 g1116(.a(new_n1324_), .O(o_59_));
  inv1 g1117(.a(i_40_), .O(new_n1326_));
  nor2 g1118(.a(new_n885_), .b(new_n1326_), .O(new_n1327_));
  nor2 g1119(.a(new_n891_), .b(new_n599_), .O(new_n1328_));
  nor2 g1120(.a(new_n898_), .b(new_n742_), .O(new_n1329_));
  nor2 g1121(.a(new_n1329_), .b(new_n1328_), .O(new_n1330_));
  inv1 g1122(.a(new_n1330_), .O(new_n1331_));
  nor2 g1123(.a(new_n916_), .b(new_n1321_), .O(new_n1332_));
  nor2 g1124(.a(new_n904_), .b(new_n839_), .O(new_n1333_));
  nor2 g1125(.a(new_n1333_), .b(new_n1332_), .O(new_n1334_));
  inv1 g1126(.a(new_n1334_), .O(new_n1335_));
  nor2 g1127(.a(new_n1335_), .b(new_n1331_), .O(new_n1336_));
  inv1 g1128(.a(new_n1336_), .O(new_n1337_));
  nor2 g1129(.a(new_n1058_), .b(new_n692_), .O(new_n1338_));
  inv1 g1130(.a(i_96_), .O(new_n1339_));
  nor2 g1131(.a(new_n910_), .b(new_n1339_), .O(new_n1340_));
  nor2 g1132(.a(new_n894_), .b(new_n589_), .O(new_n1341_));
  nor2 g1133(.a(new_n1341_), .b(new_n1340_), .O(new_n1342_));
  inv1 g1134(.a(new_n1342_), .O(new_n1343_));
  nor2 g1135(.a(new_n1343_), .b(new_n1338_), .O(new_n1344_));
  inv1 g1136(.a(new_n1344_), .O(new_n1345_));
  nor2 g1137(.a(new_n1345_), .b(new_n1337_), .O(new_n1346_));
  inv1 g1138(.a(new_n1346_), .O(new_n1347_));
  nor2 g1139(.a(new_n1347_), .b(new_n1327_), .O(new_n1348_));
  inv1 g1140(.a(new_n1348_), .O(o_6_));
  nor2 g1141(.a(i_110_), .b(new_n301_), .O(new_n1350_));
  inv1 g1142(.a(new_n1350_), .O(new_n1351_));
  nor2 g1143(.a(new_n1351_), .b(new_n1170_), .O(new_n1352_));
  nor2 g1144(.a(new_n331_), .b(new_n303_), .O(new_n1353_));
  nor2 g1145(.a(new_n1353_), .b(new_n311_), .O(new_n1354_));
  nor2 g1146(.a(new_n1354_), .b(new_n324_), .O(new_n1355_));
  nor2 g1147(.a(new_n1355_), .b(new_n271_), .O(new_n1356_));
  nor2 g1148(.a(new_n1356_), .b(new_n316_), .O(new_n1357_));
  inv1 g1149(.a(new_n1357_), .O(new_n1358_));
  nor2 g1150(.a(new_n1358_), .b(new_n1352_), .O(new_n1359_));
  inv1 g1151(.a(new_n1359_), .O(o_81_));
  nor2 g1152(.a(new_n339_), .b(i_105_), .O(new_n1361_));
  inv1 g1153(.a(new_n1361_), .O(new_n1362_));
  nor2 g1154(.a(new_n1362_), .b(new_n787_), .O(new_n1363_));
  nor2 g1155(.a(new_n1363_), .b(new_n1282_), .O(new_n1364_));
  nor2 g1156(.a(new_n242_), .b(new_n301_), .O(new_n1365_));
  inv1 g1157(.a(new_n1365_), .O(new_n1366_));
  nor2 g1158(.a(new_n1366_), .b(new_n241_), .O(new_n1367_));
  inv1 g1159(.a(new_n1367_), .O(new_n1368_));
  nor2 g1160(.a(new_n1368_), .b(new_n273_), .O(new_n1369_));
  inv1 g1161(.a(new_n1369_), .O(new_n1370_));
  nor2 g1162(.a(new_n1370_), .b(new_n257_), .O(new_n1371_));
  inv1 g1163(.a(new_n1371_), .O(new_n1372_));
  nor2 g1164(.a(new_n1372_), .b(new_n286_), .O(new_n1373_));
  nor2 g1165(.a(new_n1373_), .b(new_n335_), .O(new_n1374_));
  nor2 g1166(.a(new_n1374_), .b(new_n316_), .O(new_n1375_));
  inv1 g1167(.a(new_n1375_), .O(new_n1376_));
  nor2 g1168(.a(new_n1376_), .b(new_n1364_), .O(new_n1377_));
  inv1 g1169(.a(new_n1377_), .O(o_76_));
  inv1 g1170(.a(i_10_), .O(new_n1379_));
  inv1 g1171(.a(new_n372_), .O(new_n1380_));
  nor2 g1172(.a(new_n1380_), .b(i_80_), .O(new_n1381_));
  nor2 g1173(.a(new_n569_), .b(i_18_), .O(new_n1382_));
  inv1 g1174(.a(new_n1382_), .O(new_n1383_));
  nor2 g1175(.a(new_n1383_), .b(new_n1305_), .O(new_n1384_));
  inv1 g1176(.a(new_n1384_), .O(new_n1385_));
  nor2 g1177(.a(new_n1385_), .b(new_n1303_), .O(new_n1386_));
  nor2 g1178(.a(new_n1386_), .b(new_n1381_), .O(new_n1387_));
  nor2 g1179(.a(new_n1387_), .b(new_n1379_), .O(new_n1388_));
  nor2 g1180(.a(new_n381_), .b(new_n365_), .O(new_n1389_));
  nor2 g1181(.a(new_n227_), .b(new_n1379_), .O(new_n1390_));
  inv1 g1182(.a(new_n1390_), .O(new_n1391_));
  nor2 g1183(.a(new_n1391_), .b(i_80_), .O(new_n1392_));
  inv1 g1184(.a(new_n1392_), .O(new_n1393_));
  nor2 g1185(.a(new_n1393_), .b(new_n1389_), .O(new_n1394_));
  nor2 g1186(.a(new_n746_), .b(new_n405_), .O(new_n1395_));
  nor2 g1187(.a(new_n428_), .b(new_n1339_), .O(new_n1396_));
  nor2 g1188(.a(new_n1396_), .b(new_n1395_), .O(new_n1397_));
  inv1 g1189(.a(new_n1397_), .O(new_n1398_));
  nor2 g1190(.a(new_n1398_), .b(new_n1394_), .O(new_n1399_));
  inv1 g1191(.a(new_n1399_), .O(new_n1400_));
  nor2 g1192(.a(new_n1400_), .b(new_n1388_), .O(new_n1401_));
  inv1 g1193(.a(new_n1401_), .O(o_67_));
  inv1 g1194(.a(i_37_), .O(new_n1403_));
  nor2 g1195(.a(new_n885_), .b(new_n1403_), .O(new_n1404_));
  nor2 g1196(.a(new_n894_), .b(new_n555_), .O(new_n1405_));
  nor2 g1197(.a(new_n904_), .b(new_n845_), .O(new_n1406_));
  nor2 g1198(.a(new_n1406_), .b(new_n1405_), .O(new_n1407_));
  inv1 g1199(.a(new_n1407_), .O(new_n1408_));
  nor2 g1200(.a(new_n916_), .b(new_n735_), .O(new_n1409_));
  nor2 g1201(.a(new_n898_), .b(new_n638_), .O(new_n1410_));
  nor2 g1202(.a(new_n1410_), .b(new_n1409_), .O(new_n1411_));
  inv1 g1203(.a(new_n1411_), .O(new_n1412_));
  nor2 g1204(.a(new_n1412_), .b(new_n1408_), .O(new_n1413_));
  inv1 g1205(.a(new_n1413_), .O(new_n1414_));
  nor2 g1206(.a(new_n1058_), .b(new_n626_), .O(new_n1415_));
  nor2 g1207(.a(new_n891_), .b(new_n673_), .O(new_n1416_));
  nor2 g1208(.a(new_n910_), .b(new_n1137_), .O(new_n1417_));
  nor2 g1209(.a(new_n1417_), .b(new_n1416_), .O(new_n1418_));
  inv1 g1210(.a(new_n1418_), .O(new_n1419_));
  nor2 g1211(.a(new_n1419_), .b(new_n1415_), .O(new_n1420_));
  inv1 g1212(.a(new_n1420_), .O(new_n1421_));
  nor2 g1213(.a(new_n1421_), .b(new_n1414_), .O(new_n1422_));
  inv1 g1214(.a(new_n1422_), .O(new_n1423_));
  nor2 g1215(.a(new_n1423_), .b(new_n1404_), .O(new_n1424_));
  inv1 g1216(.a(new_n1424_), .O(o_3_));
  nor2 g1217(.a(new_n1172_), .b(i_111_), .O(new_n1426_));
  nor2 g1218(.a(new_n1355_), .b(new_n276_), .O(new_n1427_));
  nor2 g1219(.a(new_n1427_), .b(new_n316_), .O(new_n1428_));
  inv1 g1220(.a(new_n1428_), .O(new_n1429_));
  nor2 g1221(.a(new_n1429_), .b(new_n1426_), .O(new_n1430_));
  inv1 g1222(.a(new_n1430_), .O(o_82_));
  nor2 g1223(.a(new_n257_), .b(new_n237_), .O(new_n1432_));
  nor2 g1224(.a(new_n311_), .b(new_n248_), .O(new_n1433_));
  inv1 g1225(.a(new_n1433_), .O(new_n1434_));
  nor2 g1226(.a(new_n1434_), .b(new_n1432_), .O(new_n1435_));
  nor2 g1227(.a(new_n253_), .b(i_104_), .O(new_n1436_));
  inv1 g1228(.a(new_n1436_), .O(new_n1437_));
  nor2 g1229(.a(new_n1437_), .b(new_n786_), .O(new_n1438_));
  nor2 g1230(.a(new_n1438_), .b(new_n316_), .O(new_n1439_));
  inv1 g1231(.a(new_n1439_), .O(new_n1440_));
  nor2 g1232(.a(new_n1440_), .b(new_n1435_), .O(new_n1441_));
  inv1 g1233(.a(new_n1441_), .O(o_75_));
  nor2 g1234(.a(i_11_), .b(i_89_), .O(new_n1443_));
  inv1 g1235(.a(i_11_), .O(new_n1444_));
  nor2 g1236(.a(new_n1444_), .b(new_n448_), .O(new_n1445_));
  nor2 g1237(.a(new_n1445_), .b(new_n1443_), .O(new_n1446_));
  inv1 g1238(.a(new_n1446_), .O(new_n1447_));
  nor2 g1239(.a(new_n1447_), .b(i_23_), .O(new_n1448_));
  nor2 g1240(.a(new_n376_), .b(i_81_), .O(new_n1449_));
  inv1 g1241(.a(new_n1449_), .O(new_n1450_));
  nor2 g1242(.a(new_n1450_), .b(new_n1444_), .O(new_n1451_));
  nor2 g1243(.a(new_n1451_), .b(new_n1448_), .O(new_n1452_));
  nor2 g1244(.a(new_n1452_), .b(i_19_), .O(new_n1453_));
  inv1 g1245(.a(new_n1453_), .O(new_n1454_));
  nor2 g1246(.a(new_n1454_), .b(new_n409_), .O(new_n1455_));
  nor2 g1247(.a(new_n453_), .b(i_11_), .O(new_n1456_));
  inv1 g1248(.a(new_n1456_), .O(new_n1457_));
  nor2 g1249(.a(new_n1457_), .b(new_n1450_), .O(new_n1458_));
  inv1 g1250(.a(new_n1458_), .O(new_n1459_));
  nor2 g1251(.a(new_n1459_), .b(new_n397_), .O(new_n1460_));
  inv1 g1252(.a(new_n1460_), .O(new_n1461_));
  nor2 g1253(.a(new_n1461_), .b(new_n405_), .O(new_n1462_));
  nor2 g1254(.a(new_n1462_), .b(new_n1455_), .O(new_n1463_));
  nor2 g1255(.a(new_n1463_), .b(i_33_), .O(new_n1464_));
  nor2 g1256(.a(new_n1447_), .b(i_81_), .O(new_n1465_));
  inv1 g1257(.a(new_n1465_), .O(new_n1466_));
  nor2 g1258(.a(new_n1466_), .b(new_n384_), .O(new_n1467_));
  nor2 g1259(.a(new_n428_), .b(new_n1078_), .O(new_n1468_));
  nor2 g1260(.a(new_n762_), .b(new_n405_), .O(new_n1469_));
  inv1 g1261(.a(new_n367_), .O(new_n1470_));
  nor2 g1262(.a(new_n1466_), .b(new_n1470_), .O(new_n1471_));
  nor2 g1263(.a(new_n1471_), .b(new_n1469_), .O(new_n1472_));
  inv1 g1264(.a(new_n1472_), .O(new_n1473_));
  nor2 g1265(.a(new_n1473_), .b(new_n1468_), .O(new_n1474_));
  inv1 g1266(.a(new_n1474_), .O(new_n1475_));
  nor2 g1267(.a(new_n1475_), .b(new_n1467_), .O(new_n1476_));
  inv1 g1268(.a(new_n1476_), .O(new_n1477_));
  nor2 g1269(.a(new_n1477_), .b(new_n1464_), .O(new_n1478_));
  inv1 g1270(.a(new_n1478_), .O(o_68_));
  inv1 g1271(.a(i_38_), .O(new_n1480_));
  nor2 g1272(.a(new_n885_), .b(new_n1480_), .O(new_n1481_));
  nor2 g1273(.a(new_n891_), .b(new_n655_), .O(new_n1482_));
  nor2 g1274(.a(new_n898_), .b(new_n773_), .O(new_n1483_));
  nor2 g1275(.a(new_n1483_), .b(new_n1482_), .O(new_n1484_));
  inv1 g1276(.a(new_n1484_), .O(new_n1485_));
  nor2 g1277(.a(new_n916_), .b(new_n804_), .O(new_n1486_));
  nor2 g1278(.a(new_n904_), .b(new_n1049_), .O(new_n1487_));
  nor2 g1279(.a(new_n1487_), .b(new_n1486_), .O(new_n1488_));
  inv1 g1280(.a(new_n1488_), .O(new_n1489_));
  nor2 g1281(.a(new_n1489_), .b(new_n1485_), .O(new_n1490_));
  inv1 g1282(.a(new_n1490_), .O(new_n1491_));
  nor2 g1283(.a(new_n1058_), .b(new_n663_), .O(new_n1492_));
  nor2 g1284(.a(new_n910_), .b(new_n1226_), .O(new_n1493_));
  nor2 g1285(.a(new_n894_), .b(new_n526_), .O(new_n1494_));
  nor2 g1286(.a(new_n1494_), .b(new_n1493_), .O(new_n1495_));
  inv1 g1287(.a(new_n1495_), .O(new_n1496_));
  nor2 g1288(.a(new_n1496_), .b(new_n1492_), .O(new_n1497_));
  inv1 g1289(.a(new_n1497_), .O(new_n1498_));
  nor2 g1290(.a(new_n1498_), .b(new_n1491_), .O(new_n1499_));
  inv1 g1291(.a(new_n1499_), .O(new_n1500_));
  nor2 g1292(.a(new_n1500_), .b(new_n1481_), .O(new_n1501_));
  inv1 g1293(.a(new_n1501_), .O(o_4_));
  zero g1294(.O(o_29_));
  zero g1295(.O(o_31_));
  zero g1296(.O(o_30_));
  buf  g1297(.a(i_87_), .O(o_19_));
  buf  g1298(.a(i_92_), .O(o_0_));
  buf  g1299(.a(i_88_), .O(o_20_));
endmodule


