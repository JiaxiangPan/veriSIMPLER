// Benchmark "top" written by ABC on Wed Jan 17 21:32:51 2024

module top ( 
    i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_,
    o_0_  );
  input  i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;
  output o_0_;
  wire new_n11_, new_n12_, new_n13_, new_n14_, new_n15_, new_n16_, new_n17_,
    new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_, new_n24_,
    new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_, new_n31_,
    new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_, new_n38_,
    new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_,
    new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_,
    new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_;
  inv1 g000(.a(i_5_), .O(new_n11_));
  nor2 g001(.a(i_0_), .b(new_n11_), .O(new_n12_));
  inv1 g002(.a(new_n12_), .O(new_n13_));
  inv1 g003(.a(i_8_), .O(new_n14_));
  nor2 g004(.a(new_n14_), .b(i_7_), .O(new_n15_));
  inv1 g005(.a(new_n15_), .O(new_n16_));
  inv1 g006(.a(i_3_), .O(new_n17_));
  nor2 g007(.a(i_2_), .b(new_n17_), .O(new_n18_));
  inv1 g008(.a(new_n18_), .O(new_n19_));
  nor2 g009(.a(new_n19_), .b(new_n16_), .O(new_n20_));
  inv1 g010(.a(i_2_), .O(new_n21_));
  nor2 g011(.a(new_n21_), .b(new_n17_), .O(new_n22_));
  inv1 g012(.a(new_n22_), .O(new_n23_));
  nor2 g013(.a(i_8_), .b(i_7_), .O(new_n24_));
  inv1 g014(.a(new_n24_), .O(new_n25_));
  nor2 g015(.a(new_n25_), .b(new_n23_), .O(new_n26_));
  nor2 g016(.a(new_n26_), .b(new_n20_), .O(new_n27_));
  nor2 g017(.a(new_n27_), .b(new_n13_), .O(new_n28_));
  inv1 g018(.a(i_7_), .O(new_n29_));
  nor2 g019(.a(i_1_), .b(new_n29_), .O(new_n30_));
  inv1 g020(.a(new_n30_), .O(new_n31_));
  inv1 g021(.a(i_0_), .O(new_n32_));
  nor2 g022(.a(new_n32_), .b(i_4_), .O(new_n33_));
  inv1 g023(.a(new_n33_), .O(new_n34_));
  inv1 g024(.a(i_6_), .O(new_n35_));
  nor2 g025(.a(new_n35_), .b(i_8_), .O(new_n36_));
  inv1 g026(.a(new_n36_), .O(new_n37_));
  nor2 g027(.a(new_n37_), .b(new_n34_), .O(new_n38_));
  nor2 g028(.a(i_2_), .b(new_n14_), .O(new_n39_));
  inv1 g029(.a(new_n39_), .O(new_n40_));
  nor2 g030(.a(i_4_), .b(new_n35_), .O(new_n41_));
  inv1 g031(.a(new_n41_), .O(new_n42_));
  nor2 g032(.a(new_n42_), .b(new_n40_), .O(new_n43_));
  nor2 g033(.a(new_n43_), .b(new_n38_), .O(new_n44_));
  nor2 g034(.a(new_n44_), .b(new_n31_), .O(new_n45_));
  nor2 g035(.a(new_n45_), .b(new_n28_), .O(new_n46_));
  inv1 g036(.a(new_n46_), .O(new_n47_));
  nor2 g037(.a(new_n14_), .b(new_n29_), .O(new_n48_));
  inv1 g038(.a(new_n48_), .O(new_n49_));
  nor2 g039(.a(i_1_), .b(new_n11_), .O(new_n50_));
  inv1 g040(.a(new_n50_), .O(new_n51_));
  nor2 g041(.a(i_4_), .b(i_3_), .O(new_n52_));
  inv1 g042(.a(new_n52_), .O(new_n53_));
  nor2 g043(.a(new_n53_), .b(new_n51_), .O(new_n54_));
  nor2 g044(.a(new_n17_), .b(i_5_), .O(new_n55_));
  inv1 g045(.a(new_n55_), .O(new_n56_));
  nor2 g046(.a(i_0_), .b(i_4_), .O(new_n57_));
  inv1 g047(.a(new_n57_), .O(new_n58_));
  nor2 g048(.a(new_n58_), .b(new_n56_), .O(new_n59_));
  nor2 g049(.a(new_n59_), .b(new_n54_), .O(new_n60_));
  nor2 g050(.a(new_n60_), .b(new_n49_), .O(new_n61_));
  nor2 g051(.a(new_n11_), .b(i_7_), .O(new_n62_));
  inv1 g052(.a(new_n62_), .O(new_n63_));
  nor2 g053(.a(new_n63_), .b(i_4_), .O(new_n64_));
  inv1 g054(.a(i_1_), .O(new_n65_));
  nor2 g055(.a(new_n65_), .b(i_3_), .O(new_n66_));
  inv1 g056(.a(new_n66_), .O(new_n67_));
  nor2 g057(.a(new_n67_), .b(i_0_), .O(new_n68_));
  inv1 g058(.a(new_n68_), .O(new_n69_));
  nor2 g059(.a(new_n48_), .b(new_n11_), .O(new_n70_));
  inv1 g060(.a(new_n70_), .O(new_n71_));
  nor2 g061(.a(new_n71_), .b(new_n69_), .O(new_n72_));
  inv1 g062(.a(new_n72_), .O(new_n73_));
  nor2 g063(.a(new_n73_), .b(new_n64_), .O(new_n74_));
  nor2 g064(.a(new_n74_), .b(new_n61_), .O(new_n75_));
  inv1 g065(.a(new_n75_), .O(new_n76_));
  nor2 g066(.a(new_n76_), .b(new_n47_), .O(new_n77_));
  inv1 g067(.a(new_n77_), .O(new_n78_));
  nor2 g068(.a(i_2_), .b(i_1_), .O(new_n79_));
  nor2 g069(.a(new_n32_), .b(new_n65_), .O(new_n80_));
  nor2 g070(.a(new_n80_), .b(new_n79_), .O(new_n81_));
  nor2 g071(.a(new_n81_), .b(new_n17_), .O(new_n82_));
  nor2 g072(.a(new_n21_), .b(new_n65_), .O(new_n83_));
  nor2 g073(.a(new_n83_), .b(i_3_), .O(new_n84_));
  nor2 g074(.a(new_n16_), .b(i_5_), .O(new_n85_));
  inv1 g075(.a(new_n85_), .O(new_n86_));
  nor2 g076(.a(new_n86_), .b(new_n84_), .O(new_n87_));
  inv1 g077(.a(new_n87_), .O(new_n88_));
  nor2 g078(.a(new_n88_), .b(new_n82_), .O(new_n89_));
  inv1 g079(.a(i_4_), .O(new_n90_));
  nor2 g080(.a(i_0_), .b(new_n90_), .O(new_n91_));
  inv1 g081(.a(new_n91_), .O(new_n92_));
  nor2 g082(.a(new_n21_), .b(i_1_), .O(new_n93_));
  inv1 g083(.a(new_n93_), .O(new_n94_));
  nor2 g084(.a(i_8_), .b(new_n29_), .O(new_n95_));
  inv1 g085(.a(new_n95_), .O(new_n96_));
  nor2 g086(.a(new_n96_), .b(new_n94_), .O(new_n97_));
  inv1 g087(.a(new_n97_), .O(new_n98_));
  nor2 g088(.a(new_n98_), .b(new_n92_), .O(new_n99_));
  nor2 g089(.a(i_1_), .b(new_n17_), .O(new_n100_));
  inv1 g090(.a(new_n100_), .O(new_n101_));
  nor2 g091(.a(new_n101_), .b(i_0_), .O(new_n102_));
  inv1 g092(.a(new_n102_), .O(new_n103_));
  nor2 g093(.a(new_n35_), .b(i_7_), .O(new_n104_));
  inv1 g094(.a(new_n104_), .O(new_n105_));
  nor2 g095(.a(new_n105_), .b(new_n11_), .O(new_n106_));
  inv1 g096(.a(new_n106_), .O(new_n107_));
  nor2 g097(.a(new_n107_), .b(new_n103_), .O(new_n108_));
  nor2 g098(.a(new_n108_), .b(new_n99_), .O(new_n109_));
  inv1 g099(.a(new_n109_), .O(new_n110_));
  nor2 g100(.a(new_n110_), .b(new_n89_), .O(new_n111_));
  inv1 g101(.a(new_n111_), .O(new_n112_));
  nor2 g102(.a(new_n32_), .b(i_6_), .O(new_n113_));
  inv1 g103(.a(new_n113_), .O(new_n114_));
  nor2 g104(.a(new_n65_), .b(i_4_), .O(new_n115_));
  inv1 g105(.a(new_n115_), .O(new_n116_));
  nor2 g106(.a(new_n116_), .b(new_n63_), .O(new_n117_));
  nor2 g107(.a(new_n21_), .b(i_3_), .O(new_n118_));
  inv1 g108(.a(new_n118_), .O(new_n119_));
  nor2 g109(.a(new_n119_), .b(new_n51_), .O(new_n120_));
  nor2 g110(.a(new_n120_), .b(new_n117_), .O(new_n121_));
  nor2 g111(.a(new_n121_), .b(new_n114_), .O(new_n122_));
  nor2 g112(.a(new_n90_), .b(i_6_), .O(new_n123_));
  inv1 g113(.a(new_n123_), .O(new_n124_));
  nor2 g114(.a(new_n69_), .b(new_n21_), .O(new_n125_));
  inv1 g115(.a(new_n125_), .O(new_n126_));
  nor2 g116(.a(new_n126_), .b(new_n124_), .O(new_n127_));
  nor2 g117(.a(new_n127_), .b(new_n122_), .O(new_n128_));
  inv1 g118(.a(new_n128_), .O(new_n129_));
  nor2 g119(.a(new_n129_), .b(new_n112_), .O(new_n130_));
  inv1 g120(.a(new_n130_), .O(new_n131_));
  nor2 g121(.a(new_n131_), .b(new_n78_), .O(new_n132_));
  inv1 g122(.a(new_n132_), .O(new_n133_));
  nor2 g123(.a(i_5_), .b(new_n29_), .O(new_n134_));
  inv1 g124(.a(new_n134_), .O(new_n135_));
  nor2 g125(.a(new_n135_), .b(i_4_), .O(new_n136_));
  nor2 g126(.a(new_n90_), .b(i_5_), .O(new_n137_));
  inv1 g127(.a(new_n137_), .O(new_n138_));
  nor2 g128(.a(new_n138_), .b(i_8_), .O(new_n139_));
  nor2 g129(.a(new_n139_), .b(new_n136_), .O(new_n140_));
  nor2 g130(.a(new_n67_), .b(new_n32_), .O(new_n141_));
  inv1 g131(.a(new_n141_), .O(new_n142_));
  nor2 g132(.a(new_n142_), .b(new_n140_), .O(new_n143_));
  nor2 g133(.a(new_n126_), .b(new_n42_), .O(new_n144_));
  nor2 g134(.a(new_n144_), .b(new_n143_), .O(new_n145_));
  inv1 g135(.a(new_n145_), .O(new_n146_));
  nor2 g136(.a(new_n32_), .b(i_2_), .O(new_n147_));
  inv1 g137(.a(new_n147_), .O(new_n148_));
  nor2 g138(.a(new_n11_), .b(new_n29_), .O(new_n149_));
  inv1 g139(.a(new_n149_), .O(new_n150_));
  nor2 g140(.a(new_n150_), .b(i_4_), .O(new_n151_));
  inv1 g141(.a(new_n151_), .O(new_n152_));
  nor2 g142(.a(new_n152_), .b(i_6_), .O(new_n153_));
  inv1 g143(.a(new_n153_), .O(new_n154_));
  nor2 g144(.a(new_n154_), .b(new_n148_), .O(new_n155_));
  nor2 g145(.a(new_n90_), .b(i_3_), .O(new_n156_));
  inv1 g146(.a(new_n156_), .O(new_n157_));
  nor2 g147(.a(new_n157_), .b(new_n21_), .O(new_n158_));
  inv1 g148(.a(new_n158_), .O(new_n159_));
  nor2 g149(.a(new_n11_), .b(i_8_), .O(new_n160_));
  inv1 g150(.a(new_n160_), .O(new_n161_));
  nor2 g151(.a(new_n161_), .b(i_6_), .O(new_n162_));
  nor2 g152(.a(new_n105_), .b(i_8_), .O(new_n163_));
  nor2 g153(.a(new_n163_), .b(new_n162_), .O(new_n164_));
  nor2 g154(.a(new_n164_), .b(new_n159_), .O(new_n165_));
  nor2 g155(.a(new_n165_), .b(new_n155_), .O(new_n166_));
  inv1 g156(.a(new_n166_), .O(new_n167_));
  nor2 g157(.a(new_n167_), .b(new_n146_), .O(new_n168_));
  inv1 g158(.a(new_n168_), .O(new_n169_));
  nor2 g159(.a(new_n154_), .b(new_n94_), .O(new_n170_));
  nor2 g160(.a(new_n101_), .b(new_n32_), .O(new_n171_));
  inv1 g161(.a(new_n171_), .O(new_n172_));
  nor2 g162(.a(new_n105_), .b(i_5_), .O(new_n173_));
  nor2 g163(.a(new_n173_), .b(new_n64_), .O(new_n174_));
  nor2 g164(.a(new_n174_), .b(new_n172_), .O(new_n175_));
  nor2 g165(.a(new_n175_), .b(new_n170_), .O(new_n176_));
  inv1 g166(.a(new_n176_), .O(new_n177_));
  nor2 g167(.a(new_n96_), .b(i_6_), .O(new_n178_));
  inv1 g168(.a(new_n178_), .O(new_n179_));
  nor2 g169(.a(new_n92_), .b(new_n17_), .O(new_n180_));
  nor2 g170(.a(new_n65_), .b(i_5_), .O(new_n181_));
  inv1 g171(.a(new_n181_), .O(new_n182_));
  nor2 g172(.a(new_n182_), .b(new_n21_), .O(new_n183_));
  nor2 g173(.a(new_n183_), .b(new_n180_), .O(new_n184_));
  nor2 g174(.a(new_n184_), .b(new_n179_), .O(new_n185_));
  nor2 g175(.a(new_n91_), .b(new_n33_), .O(new_n186_));
  nor2 g176(.a(new_n56_), .b(i_7_), .O(new_n187_));
  inv1 g177(.a(new_n187_), .O(new_n188_));
  nor2 g178(.a(new_n188_), .b(new_n65_), .O(new_n189_));
  inv1 g179(.a(new_n189_), .O(new_n190_));
  nor2 g180(.a(new_n190_), .b(new_n186_), .O(new_n191_));
  nor2 g181(.a(new_n191_), .b(new_n185_), .O(new_n192_));
  inv1 g182(.a(new_n192_), .O(new_n193_));
  nor2 g183(.a(new_n193_), .b(new_n177_), .O(new_n194_));
  inv1 g184(.a(new_n194_), .O(new_n195_));
  nor2 g185(.a(new_n195_), .b(new_n169_), .O(new_n196_));
  inv1 g186(.a(new_n196_), .O(new_n197_));
  nor2 g187(.a(new_n197_), .b(new_n133_), .O(new_n198_));
  inv1 g188(.a(new_n198_), .O(new_n199_));
  nor2 g189(.a(new_n67_), .b(new_n40_), .O(new_n200_));
  inv1 g190(.a(new_n200_), .O(new_n201_));
  nor2 g191(.a(i_0_), .b(new_n35_), .O(new_n202_));
  inv1 g192(.a(new_n202_), .O(new_n203_));
  nor2 g193(.a(new_n203_), .b(new_n201_), .O(new_n204_));
  inv1 g194(.a(new_n20_), .O(new_n205_));
  nor2 g195(.a(new_n34_), .b(new_n205_), .O(new_n206_));
  nor2 g196(.a(new_n206_), .b(new_n204_), .O(new_n207_));
  inv1 g197(.a(new_n207_), .O(new_n208_));
  nor2 g198(.a(new_n23_), .b(i_0_), .O(new_n209_));
  inv1 g199(.a(new_n209_), .O(new_n210_));
  nor2 g200(.a(new_n96_), .b(i_5_), .O(new_n211_));
  inv1 g201(.a(new_n211_), .O(new_n212_));
  nor2 g202(.a(new_n212_), .b(new_n210_), .O(new_n213_));
  nor2 g203(.a(new_n124_), .b(new_n16_), .O(new_n214_));
  inv1 g204(.a(new_n214_), .O(new_n215_));
  nor2 g205(.a(new_n215_), .b(new_n101_), .O(new_n216_));
  nor2 g206(.a(new_n216_), .b(new_n213_), .O(new_n217_));
  inv1 g207(.a(new_n217_), .O(new_n218_));
  nor2 g208(.a(new_n218_), .b(new_n208_), .O(new_n219_));
  inv1 g209(.a(new_n219_), .O(new_n220_));
  nor2 g210(.a(new_n16_), .b(new_n35_), .O(new_n221_));
  inv1 g211(.a(new_n221_), .O(new_n222_));
  nor2 g212(.a(new_n19_), .b(i_1_), .O(new_n223_));
  inv1 g213(.a(new_n223_), .O(new_n224_));
  nor2 g214(.a(new_n224_), .b(new_n222_), .O(new_n225_));
  nor2 g215(.a(new_n101_), .b(new_n37_), .O(new_n226_));
  inv1 g216(.a(new_n226_), .O(new_n227_));
  nor2 g217(.a(new_n227_), .b(new_n138_), .O(new_n228_));
  nor2 g218(.a(new_n228_), .b(new_n225_), .O(new_n229_));
  inv1 g219(.a(new_n229_), .O(new_n230_));
  nor2 g220(.a(new_n53_), .b(new_n32_), .O(new_n231_));
  inv1 g221(.a(new_n231_), .O(new_n232_));
  nor2 g222(.a(i_6_), .b(new_n14_), .O(new_n233_));
  inv1 g223(.a(new_n233_), .O(new_n234_));
  nor2 g224(.a(new_n234_), .b(new_n11_), .O(new_n235_));
  inv1 g225(.a(new_n235_), .O(new_n236_));
  nor2 g226(.a(new_n236_), .b(new_n232_), .O(new_n237_));
  nor2 g227(.a(i_2_), .b(new_n65_), .O(new_n238_));
  inv1 g228(.a(new_n238_), .O(new_n239_));
  nor2 g229(.a(new_n239_), .b(new_n138_), .O(new_n240_));
  inv1 g230(.a(new_n240_), .O(new_n241_));
  nor2 g231(.a(new_n241_), .b(new_n203_), .O(new_n242_));
  nor2 g232(.a(new_n242_), .b(new_n237_), .O(new_n243_));
  inv1 g233(.a(new_n243_), .O(new_n244_));
  nor2 g234(.a(new_n244_), .b(new_n230_), .O(new_n245_));
  inv1 g235(.a(new_n245_), .O(new_n246_));
  nor2 g236(.a(new_n246_), .b(new_n220_), .O(new_n247_));
  inv1 g237(.a(new_n247_), .O(new_n248_));
  inv1 g238(.a(new_n43_), .O(new_n249_));
  nor2 g239(.a(new_n32_), .b(i_5_), .O(new_n250_));
  nor2 g240(.a(new_n250_), .b(new_n12_), .O(new_n251_));
  nor2 g241(.a(new_n251_), .b(new_n249_), .O(new_n252_));
  nor2 g242(.a(new_n96_), .b(new_n35_), .O(new_n253_));
  inv1 g243(.a(new_n253_), .O(new_n254_));
  nor2 g244(.a(new_n182_), .b(i_2_), .O(new_n255_));
  inv1 g245(.a(new_n255_), .O(new_n256_));
  nor2 g246(.a(new_n256_), .b(new_n254_), .O(new_n257_));
  nor2 g247(.a(new_n257_), .b(new_n252_), .O(new_n258_));
  inv1 g248(.a(new_n258_), .O(new_n259_));
  nor2 g249(.a(new_n49_), .b(i_6_), .O(new_n260_));
  inv1 g250(.a(new_n260_), .O(new_n261_));
  nor2 g251(.a(new_n138_), .b(i_1_), .O(new_n262_));
  inv1 g252(.a(new_n262_), .O(new_n263_));
  nor2 g253(.a(new_n263_), .b(new_n261_), .O(new_n264_));
  nor2 g254(.a(new_n32_), .b(i_7_), .O(new_n265_));
  inv1 g255(.a(new_n265_), .O(new_n266_));
  nor2 g256(.a(new_n266_), .b(new_n124_), .O(new_n267_));
  inv1 g257(.a(new_n267_), .O(new_n268_));
  nor2 g258(.a(new_n268_), .b(new_n40_), .O(new_n269_));
  nor2 g259(.a(new_n269_), .b(new_n264_), .O(new_n270_));
  inv1 g260(.a(new_n270_), .O(new_n271_));
  nor2 g261(.a(new_n271_), .b(new_n259_), .O(new_n272_));
  inv1 g262(.a(new_n272_), .O(new_n273_));
  nor2 g263(.a(new_n157_), .b(new_n37_), .O(new_n274_));
  inv1 g264(.a(new_n274_), .O(new_n275_));
  nor2 g265(.a(new_n275_), .b(new_n148_), .O(new_n276_));
  nor2 g266(.a(new_n157_), .b(i_2_), .O(new_n277_));
  inv1 g267(.a(new_n277_), .O(new_n278_));
  nor2 g268(.a(new_n278_), .b(new_n222_), .O(new_n279_));
  nor2 g269(.a(new_n279_), .b(new_n276_), .O(new_n280_));
  inv1 g270(.a(new_n280_), .O(new_n281_));
  nor2 g271(.a(new_n232_), .b(new_n107_), .O(new_n282_));
  inv1 g272(.a(new_n26_), .O(new_n283_));
  nor2 g273(.a(new_n34_), .b(new_n283_), .O(new_n284_));
  nor2 g274(.a(new_n284_), .b(new_n282_), .O(new_n285_));
  inv1 g275(.a(new_n285_), .O(new_n286_));
  nor2 g276(.a(new_n286_), .b(new_n281_), .O(new_n287_));
  inv1 g277(.a(new_n287_), .O(new_n288_));
  nor2 g278(.a(new_n288_), .b(new_n273_), .O(new_n289_));
  inv1 g279(.a(new_n289_), .O(new_n290_));
  nor2 g280(.a(new_n290_), .b(new_n248_), .O(new_n291_));
  inv1 g281(.a(new_n291_), .O(new_n292_));
  nor2 g282(.a(new_n19_), .b(new_n65_), .O(new_n293_));
  inv1 g283(.a(new_n293_), .O(new_n294_));
  nor2 g284(.a(new_n294_), .b(new_n179_), .O(new_n295_));
  inv1 g285(.a(new_n79_), .O(new_n296_));
  inv1 g286(.a(new_n250_), .O(new_n297_));
  nor2 g287(.a(new_n297_), .b(new_n296_), .O(new_n298_));
  inv1 g288(.a(new_n298_), .O(new_n299_));
  nor2 g289(.a(new_n299_), .b(new_n49_), .O(new_n300_));
  nor2 g290(.a(new_n300_), .b(new_n295_), .O(new_n301_));
  inv1 g291(.a(new_n301_), .O(new_n302_));
  nor2 g292(.a(new_n275_), .b(new_n51_), .O(new_n303_));
  nor2 g293(.a(new_n119_), .b(i_1_), .O(new_n304_));
  inv1 g294(.a(new_n304_), .O(new_n305_));
  nor2 g295(.a(new_n35_), .b(new_n29_), .O(new_n306_));
  inv1 g296(.a(new_n306_), .O(new_n307_));
  nor2 g297(.a(new_n307_), .b(i_5_), .O(new_n308_));
  inv1 g298(.a(new_n308_), .O(new_n309_));
  nor2 g299(.a(new_n309_), .b(new_n305_), .O(new_n310_));
  nor2 g300(.a(new_n310_), .b(new_n303_), .O(new_n311_));
  inv1 g301(.a(new_n311_), .O(new_n312_));
  nor2 g302(.a(new_n312_), .b(new_n302_), .O(new_n313_));
  inv1 g303(.a(new_n313_), .O(new_n314_));
  inv1 g304(.a(new_n83_), .O(new_n315_));
  nor2 g305(.a(new_n315_), .b(i_8_), .O(new_n316_));
  inv1 g306(.a(new_n316_), .O(new_n317_));
  nor2 g307(.a(new_n317_), .b(new_n188_), .O(new_n318_));
  nor2 g308(.a(new_n116_), .b(new_n13_), .O(new_n319_));
  inv1 g309(.a(new_n319_), .O(new_n320_));
  nor2 g310(.a(new_n320_), .b(new_n234_), .O(new_n321_));
  nor2 g311(.a(new_n321_), .b(new_n318_), .O(new_n322_));
  inv1 g312(.a(new_n322_), .O(new_n323_));
  nor2 g313(.a(new_n305_), .b(new_n222_), .O(new_n324_));
  nor2 g314(.a(new_n297_), .b(new_n201_), .O(new_n325_));
  nor2 g315(.a(new_n325_), .b(new_n324_), .O(new_n326_));
  inv1 g316(.a(new_n326_), .O(new_n327_));
  nor2 g317(.a(new_n327_), .b(new_n323_), .O(new_n328_));
  inv1 g318(.a(new_n328_), .O(new_n329_));
  nor2 g319(.a(new_n329_), .b(new_n314_), .O(new_n330_));
  inv1 g320(.a(new_n330_), .O(new_n331_));
  nor2 g321(.a(new_n239_), .b(new_n67_), .O(new_n332_));
  inv1 g322(.a(new_n332_), .O(new_n333_));
  nor2 g323(.a(new_n124_), .b(new_n11_), .O(new_n334_));
  inv1 g324(.a(new_n334_), .O(new_n335_));
  nor2 g325(.a(new_n335_), .b(new_n333_), .O(new_n336_));
  nor2 g326(.a(new_n21_), .b(i_8_), .O(new_n337_));
  inv1 g327(.a(new_n337_), .O(new_n338_));
  nor2 g328(.a(new_n338_), .b(new_n268_), .O(new_n339_));
  nor2 g329(.a(new_n339_), .b(new_n336_), .O(new_n340_));
  inv1 g330(.a(new_n340_), .O(new_n341_));
  nor2 g331(.a(new_n16_), .b(i_6_), .O(new_n342_));
  inv1 g332(.a(new_n342_), .O(new_n343_));
  nor2 g333(.a(new_n343_), .b(new_n159_), .O(new_n344_));
  nor2 g334(.a(new_n234_), .b(new_n182_), .O(new_n345_));
  inv1 g335(.a(new_n345_), .O(new_n346_));
  nor2 g336(.a(new_n346_), .b(new_n119_), .O(new_n347_));
  nor2 g337(.a(new_n347_), .b(new_n344_), .O(new_n348_));
  inv1 g338(.a(new_n348_), .O(new_n349_));
  nor2 g339(.a(new_n349_), .b(new_n341_), .O(new_n350_));
  inv1 g340(.a(new_n350_), .O(new_n351_));
  nor2 g341(.a(new_n333_), .b(new_n152_), .O(new_n352_));
  inv1 g342(.a(new_n162_), .O(new_n353_));
  nor2 g343(.a(new_n116_), .b(new_n21_), .O(new_n354_));
  inv1 g344(.a(new_n354_), .O(new_n355_));
  nor2 g345(.a(new_n355_), .b(new_n353_), .O(new_n356_));
  nor2 g346(.a(new_n356_), .b(new_n352_), .O(new_n357_));
  inv1 g347(.a(new_n357_), .O(new_n358_));
  nor2 g348(.a(new_n114_), .b(new_n98_), .O(new_n359_));
  nor2 g349(.a(new_n317_), .b(new_n232_), .O(new_n360_));
  nor2 g350(.a(new_n360_), .b(new_n359_), .O(new_n361_));
  inv1 g351(.a(new_n361_), .O(new_n362_));
  nor2 g352(.a(new_n362_), .b(new_n358_), .O(new_n363_));
  inv1 g353(.a(new_n363_), .O(new_n364_));
  nor2 g354(.a(new_n364_), .b(new_n351_), .O(new_n365_));
  inv1 g355(.a(new_n365_), .O(new_n366_));
  nor2 g356(.a(new_n366_), .b(new_n331_), .O(new_n367_));
  inv1 g357(.a(new_n367_), .O(new_n368_));
  nor2 g358(.a(new_n368_), .b(new_n292_), .O(new_n369_));
  inv1 g359(.a(new_n369_), .O(new_n370_));
  nor2 g360(.a(new_n343_), .b(new_n13_), .O(new_n371_));
  inv1 g361(.a(new_n38_), .O(new_n372_));
  nor2 g362(.a(new_n372_), .b(i_5_), .O(new_n373_));
  nor2 g363(.a(new_n373_), .b(new_n371_), .O(new_n374_));
  nor2 g364(.a(new_n374_), .b(new_n21_), .O(new_n375_));
  nor2 g365(.a(new_n210_), .b(i_7_), .O(new_n376_));
  nor2 g366(.a(new_n148_), .b(new_n31_), .O(new_n377_));
  nor2 g367(.a(new_n377_), .b(new_n376_), .O(new_n378_));
  nor2 g368(.a(new_n378_), .b(new_n124_), .O(new_n379_));
  nor2 g369(.a(new_n379_), .b(new_n375_), .O(new_n380_));
  inv1 g370(.a(new_n380_), .O(new_n381_));
  nor2 g371(.a(new_n261_), .b(new_n94_), .O(new_n382_));
  inv1 g372(.a(new_n117_), .O(new_n383_));
  nor2 g373(.a(new_n383_), .b(new_n17_), .O(new_n384_));
  nor2 g374(.a(new_n384_), .b(new_n382_), .O(new_n385_));
  nor2 g375(.a(new_n385_), .b(i_0_), .O(new_n386_));
  nor2 g376(.a(new_n21_), .b(i_4_), .O(new_n387_));
  nor2 g377(.a(new_n387_), .b(new_n238_), .O(new_n388_));
  nor2 g378(.a(new_n388_), .b(new_n37_), .O(new_n389_));
  nor2 g379(.a(new_n157_), .b(new_n31_), .O(new_n390_));
  nor2 g380(.a(new_n390_), .b(new_n389_), .O(new_n391_));
  nor2 g381(.a(new_n391_), .b(new_n13_), .O(new_n392_));
  nor2 g382(.a(new_n392_), .b(new_n386_), .O(new_n393_));
  inv1 g383(.a(new_n393_), .O(new_n394_));
  nor2 g384(.a(new_n394_), .b(new_n381_), .O(new_n395_));
  inv1 g385(.a(new_n395_), .O(new_n396_));
  nor2 g386(.a(new_n92_), .b(i_2_), .O(new_n397_));
  inv1 g387(.a(new_n397_), .O(new_n398_));
  nor2 g388(.a(new_n398_), .b(new_n236_), .O(new_n399_));
  nor2 g389(.a(new_n92_), .b(new_n296_), .O(new_n400_));
  inv1 g390(.a(new_n400_), .O(new_n401_));
  nor2 g391(.a(new_n401_), .b(new_n307_), .O(new_n402_));
  nor2 g392(.a(new_n402_), .b(new_n399_), .O(new_n403_));
  inv1 g393(.a(new_n403_), .O(new_n404_));
  nor2 g394(.a(new_n138_), .b(new_n29_), .O(new_n405_));
  inv1 g395(.a(new_n405_), .O(new_n406_));
  nor2 g396(.a(new_n406_), .b(new_n69_), .O(new_n407_));
  nor2 g397(.a(new_n296_), .b(new_n11_), .O(new_n408_));
  inv1 g398(.a(new_n408_), .O(new_n409_));
  nor2 g399(.a(new_n157_), .b(new_n32_), .O(new_n410_));
  inv1 g400(.a(new_n410_), .O(new_n411_));
  nor2 g401(.a(new_n411_), .b(new_n409_), .O(new_n412_));
  nor2 g402(.a(new_n412_), .b(new_n407_), .O(new_n413_));
  inv1 g403(.a(new_n413_), .O(new_n414_));
  nor2 g404(.a(new_n414_), .b(new_n404_), .O(new_n415_));
  inv1 g405(.a(new_n415_), .O(new_n416_));
  nor2 g406(.a(new_n309_), .b(new_n103_), .O(new_n417_));
  nor2 g407(.a(new_n90_), .b(new_n11_), .O(new_n418_));
  inv1 g408(.a(new_n418_), .O(new_n419_));
  nor2 g409(.a(new_n419_), .b(new_n19_), .O(new_n420_));
  inv1 g410(.a(new_n420_), .O(new_n421_));
  nor2 g411(.a(new_n421_), .b(new_n25_), .O(new_n422_));
  nor2 g412(.a(new_n422_), .b(new_n417_), .O(new_n423_));
  inv1 g413(.a(new_n423_), .O(new_n424_));
  nor2 g414(.a(new_n261_), .b(new_n256_), .O(new_n425_));
  nor2 g415(.a(new_n346_), .b(new_n92_), .O(new_n426_));
  nor2 g416(.a(new_n426_), .b(new_n425_), .O(new_n427_));
  inv1 g417(.a(new_n427_), .O(new_n428_));
  nor2 g418(.a(new_n428_), .b(new_n424_), .O(new_n429_));
  inv1 g419(.a(new_n429_), .O(new_n430_));
  nor2 g420(.a(new_n430_), .b(new_n416_), .O(new_n431_));
  inv1 g421(.a(new_n431_), .O(new_n432_));
  inv1 g422(.a(new_n173_), .O(new_n433_));
  nor2 g423(.a(new_n294_), .b(new_n433_), .O(new_n434_));
  nor2 g424(.a(new_n268_), .b(new_n56_), .O(new_n435_));
  nor2 g425(.a(new_n435_), .b(new_n434_), .O(new_n436_));
  inv1 g426(.a(new_n436_), .O(new_n437_));
  nor2 g427(.a(new_n239_), .b(new_n372_), .O(new_n438_));
  nor2 g428(.a(i_1_), .b(new_n35_), .O(new_n439_));
  inv1 g429(.a(new_n439_), .O(new_n440_));
  nor2 g430(.a(new_n440_), .b(new_n283_), .O(new_n441_));
  nor2 g431(.a(new_n441_), .b(new_n438_), .O(new_n442_));
  inv1 g432(.a(new_n442_), .O(new_n443_));
  nor2 g433(.a(new_n443_), .b(new_n437_), .O(new_n444_));
  inv1 g434(.a(new_n444_), .O(new_n445_));
  nor2 g435(.a(new_n409_), .b(new_n254_), .O(new_n446_));
  inv1 g436(.a(new_n387_), .O(new_n447_));
  nor2 g437(.a(new_n297_), .b(new_n234_), .O(new_n448_));
  inv1 g438(.a(new_n448_), .O(new_n449_));
  nor2 g439(.a(new_n449_), .b(new_n447_), .O(new_n450_));
  nor2 g440(.a(new_n450_), .b(new_n446_), .O(new_n451_));
  inv1 g441(.a(new_n451_), .O(new_n452_));
  inv1 g442(.a(new_n136_), .O(new_n453_));
  nor2 g443(.a(new_n172_), .b(new_n453_), .O(new_n454_));
  nor2 g444(.a(new_n152_), .b(new_n103_), .O(new_n455_));
  nor2 g445(.a(new_n455_), .b(new_n454_), .O(new_n456_));
  inv1 g446(.a(new_n456_), .O(new_n457_));
  nor2 g447(.a(new_n457_), .b(new_n452_), .O(new_n458_));
  inv1 g448(.a(new_n458_), .O(new_n459_));
  nor2 g449(.a(new_n459_), .b(new_n445_), .O(new_n460_));
  inv1 g450(.a(new_n460_), .O(new_n461_));
  nor2 g451(.a(new_n461_), .b(new_n432_), .O(new_n462_));
  inv1 g452(.a(new_n462_), .O(new_n463_));
  nor2 g453(.a(new_n463_), .b(new_n396_), .O(new_n464_));
  inv1 g454(.a(new_n464_), .O(new_n465_));
  nor2 g455(.a(new_n465_), .b(new_n370_), .O(new_n466_));
  inv1 g456(.a(new_n466_), .O(new_n467_));
  nor2 g457(.a(new_n467_), .b(new_n199_), .O(new_n468_));
  inv1 g458(.a(new_n468_), .O(o_0_));
endmodule


