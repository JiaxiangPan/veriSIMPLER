// Benchmark "top" written by ABC on Wed Jan 17 21:32:49 2024

module top ( 
    i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_,
    o_1_, o_2_, o_0_, o_3_  );
  input  i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;
  output o_1_, o_2_, o_0_, o_3_;
  wire new_n15_, new_n16_, new_n17_, new_n18_, new_n19_, new_n20_, new_n21_,
    new_n22_, new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_,
    new_n29_, new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_,
    new_n36_, new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_,
    new_n43_, new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_,
    new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_;
  inv1 g000(.a(i_0_), .O(new_n15_));
  nor2 g001(.a(new_n15_), .b(i_9_), .O(new_n16_));
  inv1 g002(.a(new_n16_), .O(new_n17_));
  inv1 g003(.a(i_2_), .O(new_n18_));
  nor2 g004(.a(new_n18_), .b(i_1_), .O(new_n19_));
  inv1 g005(.a(new_n19_), .O(new_n20_));
  nor2 g006(.a(new_n20_), .b(new_n17_), .O(new_n21_));
  inv1 g007(.a(new_n21_), .O(new_n22_));
  inv1 g008(.a(i_6_), .O(new_n23_));
  inv1 g009(.a(i_7_), .O(new_n24_));
  inv1 g010(.a(i_8_), .O(new_n25_));
  nor2 g011(.a(new_n25_), .b(new_n24_), .O(new_n26_));
  inv1 g012(.a(new_n26_), .O(new_n27_));
  nor2 g013(.a(new_n27_), .b(new_n23_), .O(new_n28_));
  inv1 g014(.a(new_n28_), .O(new_n29_));
  inv1 g015(.a(i_3_), .O(new_n30_));
  inv1 g016(.a(i_4_), .O(new_n31_));
  nor2 g017(.a(new_n31_), .b(i_5_), .O(new_n32_));
  inv1 g018(.a(new_n32_), .O(new_n33_));
  nor2 g019(.a(new_n33_), .b(new_n30_), .O(new_n34_));
  inv1 g020(.a(new_n34_), .O(new_n35_));
  nor2 g021(.a(new_n35_), .b(new_n29_), .O(new_n36_));
  nor2 g022(.a(i_8_), .b(new_n24_), .O(new_n37_));
  inv1 g023(.a(new_n37_), .O(new_n38_));
  nor2 g024(.a(new_n38_), .b(i_6_), .O(new_n39_));
  inv1 g025(.a(new_n39_), .O(new_n40_));
  nor2 g026(.a(i_3_), .b(i_5_), .O(new_n41_));
  inv1 g027(.a(new_n41_), .O(new_n42_));
  nor2 g028(.a(new_n42_), .b(i_4_), .O(new_n43_));
  inv1 g029(.a(new_n43_), .O(new_n44_));
  nor2 g030(.a(new_n44_), .b(new_n40_), .O(new_n45_));
  nor2 g031(.a(new_n45_), .b(new_n36_), .O(new_n46_));
  nor2 g032(.a(new_n46_), .b(new_n22_), .O(new_n47_));
  nor2 g033(.a(new_n30_), .b(i_5_), .O(new_n48_));
  inv1 g034(.a(new_n48_), .O(new_n49_));
  nor2 g035(.a(new_n49_), .b(i_4_), .O(new_n50_));
  inv1 g036(.a(new_n50_), .O(new_n51_));
  nor2 g037(.a(i_8_), .b(i_9_), .O(new_n52_));
  inv1 g038(.a(new_n52_), .O(new_n53_));
  nor2 g039(.a(new_n53_), .b(i_0_), .O(new_n54_));
  inv1 g040(.a(new_n54_), .O(new_n55_));
  nor2 g041(.a(i_2_), .b(i_1_), .O(new_n56_));
  inv1 g042(.a(new_n56_), .O(new_n57_));
  nor2 g043(.a(new_n57_), .b(i_6_), .O(new_n58_));
  inv1 g044(.a(new_n58_), .O(new_n59_));
  nor2 g045(.a(new_n59_), .b(new_n55_), .O(new_n60_));
  inv1 g046(.a(new_n60_), .O(new_n61_));
  nor2 g047(.a(new_n61_), .b(new_n51_), .O(new_n62_));
  inv1 g048(.a(new_n62_), .O(new_n63_));
  nor2 g049(.a(new_n63_), .b(i_7_), .O(new_n64_));
  inv1 g050(.a(i_1_), .O(new_n65_));
  nor2 g051(.a(new_n18_), .b(new_n65_), .O(new_n66_));
  inv1 g052(.a(new_n66_), .O(new_n67_));
  nor2 g053(.a(new_n67_), .b(new_n17_), .O(new_n68_));
  inv1 g054(.a(new_n68_), .O(new_n69_));
  nor2 g055(.a(new_n51_), .b(new_n29_), .O(new_n70_));
  nor2 g056(.a(new_n27_), .b(i_6_), .O(new_n71_));
  inv1 g057(.a(new_n71_), .O(new_n72_));
  nor2 g058(.a(new_n72_), .b(new_n35_), .O(new_n73_));
  nor2 g059(.a(new_n73_), .b(new_n70_), .O(new_n74_));
  nor2 g060(.a(new_n74_), .b(new_n69_), .O(new_n75_));
  nor2 g061(.a(new_n75_), .b(new_n64_), .O(new_n76_));
  inv1 g062(.a(new_n76_), .O(new_n77_));
  nor2 g063(.a(new_n77_), .b(new_n47_), .O(new_n78_));
  inv1 g064(.a(new_n78_), .O(new_n79_));
  inv1 g065(.a(new_n36_), .O(new_n80_));
  nor2 g066(.a(i_2_), .b(new_n65_), .O(new_n81_));
  inv1 g067(.a(new_n81_), .O(new_n82_));
  nor2 g068(.a(new_n82_), .b(new_n17_), .O(new_n83_));
  inv1 g069(.a(new_n83_), .O(new_n84_));
  nor2 g070(.a(new_n84_), .b(new_n80_), .O(new_n85_));
  inv1 g071(.a(new_n45_), .O(new_n86_));
  nor2 g072(.a(new_n61_), .b(new_n86_), .O(new_n87_));
  nor2 g073(.a(new_n87_), .b(new_n85_), .O(new_n88_));
  inv1 g074(.a(new_n88_), .O(new_n89_));
  nor2 g075(.a(new_n51_), .b(new_n40_), .O(new_n90_));
  inv1 g076(.a(new_n90_), .O(new_n91_));
  nor2 g077(.a(new_n82_), .b(i_9_), .O(new_n92_));
  inv1 g078(.a(new_n92_), .O(new_n93_));
  nor2 g079(.a(new_n93_), .b(i_0_), .O(new_n94_));
  inv1 g080(.a(new_n94_), .O(new_n95_));
  nor2 g081(.a(new_n95_), .b(new_n91_), .O(new_n96_));
  nor2 g082(.a(new_n82_), .b(i_0_), .O(new_n97_));
  inv1 g083(.a(new_n97_), .O(new_n98_));
  nor2 g084(.a(new_n25_), .b(i_7_), .O(new_n99_));
  inv1 g085(.a(new_n99_), .O(new_n100_));
  nor2 g086(.a(i_6_), .b(i_9_), .O(new_n101_));
  inv1 g087(.a(new_n101_), .O(new_n102_));
  nor2 g088(.a(new_n102_), .b(new_n100_), .O(new_n103_));
  inv1 g089(.a(new_n103_), .O(new_n104_));
  nor2 g090(.a(new_n104_), .b(new_n51_), .O(new_n105_));
  inv1 g091(.a(new_n105_), .O(new_n106_));
  nor2 g092(.a(new_n106_), .b(new_n98_), .O(new_n107_));
  nor2 g093(.a(new_n107_), .b(new_n96_), .O(new_n108_));
  inv1 g094(.a(new_n108_), .O(new_n109_));
  nor2 g095(.a(new_n109_), .b(new_n89_), .O(new_n110_));
  inv1 g096(.a(new_n110_), .O(new_n111_));
  nor2 g097(.a(new_n57_), .b(new_n17_), .O(new_n112_));
  inv1 g098(.a(new_n112_), .O(new_n113_));
  nor2 g099(.a(new_n113_), .b(new_n91_), .O(new_n114_));
  nor2 g100(.a(new_n33_), .b(i_3_), .O(new_n115_));
  inv1 g101(.a(new_n115_), .O(new_n116_));
  nor2 g102(.a(new_n69_), .b(new_n29_), .O(new_n117_));
  inv1 g103(.a(new_n117_), .O(new_n118_));
  nor2 g104(.a(new_n118_), .b(new_n116_), .O(new_n119_));
  nor2 g105(.a(new_n119_), .b(new_n114_), .O(new_n120_));
  inv1 g106(.a(new_n120_), .O(new_n121_));
  nor2 g107(.a(new_n38_), .b(new_n23_), .O(new_n122_));
  inv1 g108(.a(new_n122_), .O(new_n123_));
  nor2 g109(.a(new_n116_), .b(new_n22_), .O(new_n124_));
  inv1 g110(.a(new_n124_), .O(new_n125_));
  nor2 g111(.a(new_n125_), .b(new_n123_), .O(new_n126_));
  nor2 g112(.a(new_n100_), .b(new_n23_), .O(new_n127_));
  inv1 g113(.a(new_n127_), .O(new_n128_));
  nor2 g114(.a(new_n128_), .b(new_n69_), .O(new_n129_));
  inv1 g115(.a(new_n129_), .O(new_n130_));
  nor2 g116(.a(new_n130_), .b(new_n35_), .O(new_n131_));
  nor2 g117(.a(new_n131_), .b(new_n126_), .O(new_n132_));
  inv1 g118(.a(new_n132_), .O(new_n133_));
  nor2 g119(.a(new_n133_), .b(new_n121_), .O(new_n134_));
  inv1 g120(.a(new_n134_), .O(new_n135_));
  nor2 g121(.a(new_n135_), .b(new_n111_), .O(new_n136_));
  inv1 g122(.a(new_n136_), .O(new_n137_));
  nor2 g123(.a(i_0_), .b(i_9_), .O(new_n138_));
  inv1 g124(.a(new_n138_), .O(new_n139_));
  nor2 g125(.a(new_n139_), .b(new_n67_), .O(new_n140_));
  inv1 g126(.a(new_n140_), .O(new_n141_));
  nor2 g127(.a(new_n141_), .b(new_n29_), .O(new_n142_));
  nor2 g128(.a(new_n123_), .b(new_n69_), .O(new_n143_));
  nor2 g129(.a(new_n40_), .b(new_n22_), .O(new_n144_));
  nor2 g130(.a(new_n144_), .b(new_n143_), .O(new_n145_));
  inv1 g131(.a(new_n145_), .O(new_n146_));
  nor2 g132(.a(new_n146_), .b(new_n142_), .O(new_n147_));
  nor2 g133(.a(new_n147_), .b(new_n35_), .O(new_n148_));
  nor2 g134(.a(new_n91_), .b(new_n69_), .O(new_n149_));
  inv1 g135(.a(new_n70_), .O(new_n150_));
  nor2 g136(.a(new_n95_), .b(new_n150_), .O(new_n151_));
  nor2 g137(.a(new_n151_), .b(new_n149_), .O(new_n152_));
  inv1 g138(.a(new_n152_), .O(new_n153_));
  nor2 g139(.a(new_n98_), .b(new_n35_), .O(new_n154_));
  inv1 g140(.a(new_n154_), .O(new_n155_));
  nor2 g141(.a(new_n25_), .b(i_9_), .O(new_n156_));
  inv1 g142(.a(new_n156_), .O(new_n157_));
  nor2 g143(.a(new_n157_), .b(new_n23_), .O(new_n158_));
  inv1 g144(.a(new_n158_), .O(new_n159_));
  nor2 g145(.a(new_n159_), .b(i_7_), .O(new_n160_));
  inv1 g146(.a(new_n160_), .O(new_n161_));
  nor2 g147(.a(new_n161_), .b(new_n155_), .O(new_n162_));
  nor2 g148(.a(new_n84_), .b(new_n51_), .O(new_n163_));
  inv1 g149(.a(new_n163_), .O(new_n164_));
  nor2 g150(.a(new_n164_), .b(new_n72_), .O(new_n165_));
  nor2 g151(.a(new_n165_), .b(new_n162_), .O(new_n166_));
  inv1 g152(.a(new_n166_), .O(new_n167_));
  nor2 g153(.a(new_n167_), .b(new_n153_), .O(new_n168_));
  inv1 g154(.a(new_n168_), .O(new_n169_));
  nor2 g155(.a(new_n169_), .b(new_n148_), .O(new_n170_));
  inv1 g156(.a(new_n170_), .O(new_n171_));
  nor2 g157(.a(new_n171_), .b(new_n137_), .O(new_n172_));
  inv1 g158(.a(new_n172_), .O(new_n173_));
  nor2 g159(.a(new_n173_), .b(new_n79_), .O(new_n174_));
  inv1 g160(.a(new_n174_), .O(o_1_));
  nor2 g161(.a(new_n157_), .b(i_1_), .O(new_n176_));
  inv1 g162(.a(new_n176_), .O(new_n177_));
  nor2 g163(.a(new_n18_), .b(new_n23_), .O(new_n178_));
  nor2 g164(.a(new_n178_), .b(new_n177_), .O(new_n179_));
  nor2 g165(.a(i_7_), .b(i_9_), .O(new_n180_));
  inv1 g166(.a(new_n180_), .O(new_n181_));
  nor2 g167(.a(new_n18_), .b(i_4_), .O(new_n182_));
  nor2 g168(.a(new_n31_), .b(i_6_), .O(new_n183_));
  nor2 g169(.a(new_n183_), .b(new_n182_), .O(new_n184_));
  nor2 g170(.a(new_n184_), .b(new_n181_), .O(new_n185_));
  nor2 g171(.a(new_n185_), .b(new_n179_), .O(new_n186_));
  nor2 g172(.a(new_n186_), .b(i_5_), .O(new_n187_));
  nor2 g173(.a(new_n15_), .b(new_n31_), .O(new_n188_));
  nor2 g174(.a(new_n42_), .b(new_n65_), .O(new_n189_));
  inv1 g175(.a(new_n189_), .O(new_n190_));
  nor2 g176(.a(new_n190_), .b(i_9_), .O(new_n191_));
  inv1 g177(.a(new_n191_), .O(new_n192_));
  nor2 g178(.a(new_n192_), .b(new_n188_), .O(new_n193_));
  inv1 g179(.a(new_n188_), .O(new_n194_));
  nor2 g180(.a(new_n194_), .b(new_n18_), .O(new_n195_));
  nor2 g181(.a(new_n23_), .b(i_5_), .O(new_n196_));
  inv1 g182(.a(new_n196_), .O(new_n197_));
  nor2 g183(.a(new_n197_), .b(new_n53_), .O(new_n198_));
  inv1 g184(.a(new_n198_), .O(new_n199_));
  nor2 g185(.a(new_n199_), .b(new_n195_), .O(new_n200_));
  nor2 g186(.a(i_5_), .b(i_7_), .O(new_n201_));
  inv1 g187(.a(new_n201_), .O(new_n202_));
  nor2 g188(.a(new_n202_), .b(new_n177_), .O(new_n203_));
  nor2 g189(.a(new_n203_), .b(new_n200_), .O(new_n204_));
  inv1 g190(.a(new_n204_), .O(new_n205_));
  nor2 g191(.a(new_n33_), .b(i_2_), .O(new_n206_));
  inv1 g192(.a(new_n206_), .O(new_n207_));
  nor2 g193(.a(new_n207_), .b(new_n102_), .O(new_n208_));
  inv1 g194(.a(new_n182_), .O(new_n209_));
  nor2 g195(.a(new_n139_), .b(i_5_), .O(new_n210_));
  inv1 g196(.a(new_n210_), .O(new_n211_));
  nor2 g197(.a(new_n211_), .b(new_n209_), .O(new_n212_));
  nor2 g198(.a(new_n212_), .b(new_n208_), .O(new_n213_));
  inv1 g199(.a(new_n213_), .O(new_n214_));
  nor2 g200(.a(new_n214_), .b(new_n205_), .O(new_n215_));
  inv1 g201(.a(new_n215_), .O(new_n216_));
  nor2 g202(.a(new_n216_), .b(new_n193_), .O(new_n217_));
  inv1 g203(.a(new_n217_), .O(new_n218_));
  nor2 g204(.a(new_n218_), .b(new_n187_), .O(new_n219_));
  inv1 g205(.a(new_n219_), .O(new_n220_));
  nor2 g206(.a(new_n197_), .b(new_n181_), .O(new_n221_));
  nor2 g207(.a(new_n221_), .b(new_n191_), .O(new_n222_));
  nor2 g208(.a(new_n222_), .b(i_8_), .O(new_n223_));
  nor2 g209(.a(new_n202_), .b(new_n17_), .O(new_n224_));
  nor2 g210(.a(new_n224_), .b(new_n191_), .O(new_n225_));
  nor2 g211(.a(new_n225_), .b(i_2_), .O(new_n226_));
  nor2 g212(.a(new_n226_), .b(new_n223_), .O(new_n227_));
  inv1 g213(.a(new_n227_), .O(new_n228_));
  nor2 g214(.a(new_n190_), .b(i_6_), .O(new_n229_));
  nor2 g215(.a(new_n229_), .b(i_5_), .O(new_n230_));
  nor2 g216(.a(new_n230_), .b(i_9_), .O(new_n231_));
  nor2 g217(.a(new_n188_), .b(i_5_), .O(new_n232_));
  inv1 g218(.a(new_n232_), .O(new_n233_));
  nor2 g219(.a(new_n233_), .b(new_n177_), .O(new_n234_));
  nor2 g220(.a(new_n181_), .b(i_3_), .O(new_n235_));
  nor2 g221(.a(i_0_), .b(new_n31_), .O(new_n236_));
  inv1 g222(.a(new_n236_), .O(new_n237_));
  nor2 g223(.a(new_n237_), .b(new_n102_), .O(new_n238_));
  nor2 g224(.a(new_n238_), .b(new_n235_), .O(new_n239_));
  inv1 g225(.a(new_n239_), .O(new_n240_));
  nor2 g226(.a(new_n240_), .b(new_n234_), .O(new_n241_));
  inv1 g227(.a(new_n241_), .O(new_n242_));
  nor2 g228(.a(new_n242_), .b(new_n231_), .O(new_n243_));
  inv1 g229(.a(new_n243_), .O(new_n244_));
  nor2 g230(.a(new_n244_), .b(new_n228_), .O(new_n245_));
  inv1 g231(.a(new_n245_), .O(new_n246_));
  nor2 g232(.a(new_n246_), .b(new_n220_), .O(new_n247_));
  inv1 g233(.a(new_n247_), .O(o_2_));
  nor2 g234(.a(i_6_), .b(i_5_), .O(new_n249_));
  inv1 g235(.a(new_n249_), .O(new_n250_));
  nor2 g236(.a(new_n250_), .b(i_4_), .O(new_n251_));
  inv1 g237(.a(new_n251_), .O(new_n252_));
  nor2 g238(.a(new_n30_), .b(i_7_), .O(new_n253_));
  inv1 g239(.a(new_n253_), .O(new_n254_));
  nor2 g240(.a(new_n254_), .b(i_2_), .O(new_n255_));
  inv1 g241(.a(new_n255_), .O(new_n256_));
  nor2 g242(.a(new_n256_), .b(new_n55_), .O(new_n257_));
  nor2 g243(.a(new_n65_), .b(new_n30_), .O(new_n258_));
  inv1 g244(.a(new_n258_), .O(new_n259_));
  nor2 g245(.a(new_n27_), .b(new_n17_), .O(new_n260_));
  inv1 g246(.a(new_n260_), .O(new_n261_));
  nor2 g247(.a(new_n261_), .b(new_n259_), .O(new_n262_));
  nor2 g248(.a(new_n53_), .b(new_n24_), .O(new_n263_));
  inv1 g249(.a(new_n263_), .O(new_n264_));
  nor2 g250(.a(new_n57_), .b(i_3_), .O(new_n265_));
  inv1 g251(.a(new_n265_), .O(new_n266_));
  nor2 g252(.a(new_n266_), .b(new_n264_), .O(new_n267_));
  nor2 g253(.a(new_n267_), .b(new_n262_), .O(new_n268_));
  inv1 g254(.a(new_n268_), .O(new_n269_));
  nor2 g255(.a(new_n269_), .b(new_n257_), .O(new_n270_));
  nor2 g256(.a(new_n270_), .b(new_n252_), .O(new_n271_));
  nor2 g257(.a(new_n93_), .b(new_n150_), .O(new_n272_));
  nor2 g258(.a(new_n23_), .b(new_n24_), .O(new_n273_));
  inv1 g259(.a(new_n273_), .O(new_n274_));
  nor2 g260(.a(new_n274_), .b(new_n125_), .O(new_n275_));
  nor2 g261(.a(new_n275_), .b(new_n62_), .O(new_n276_));
  inv1 g262(.a(new_n276_), .O(new_n277_));
  nor2 g263(.a(new_n277_), .b(new_n272_), .O(new_n278_));
  inv1 g264(.a(new_n278_), .O(new_n279_));
  nor2 g265(.a(new_n237_), .b(new_n202_), .O(new_n280_));
  inv1 g266(.a(new_n280_), .O(new_n281_));
  nor2 g267(.a(new_n281_), .b(new_n259_), .O(new_n282_));
  nor2 g268(.a(new_n282_), .b(new_n154_), .O(new_n283_));
  nor2 g269(.a(new_n283_), .b(new_n159_), .O(new_n284_));
  nor2 g270(.a(new_n49_), .b(i_6_), .O(new_n285_));
  inv1 g271(.a(new_n285_), .O(new_n286_));
  nor2 g272(.a(new_n286_), .b(new_n67_), .O(new_n287_));
  nor2 g273(.a(new_n35_), .b(new_n20_), .O(new_n288_));
  nor2 g274(.a(new_n288_), .b(new_n287_), .O(new_n289_));
  nor2 g275(.a(new_n264_), .b(new_n15_), .O(new_n290_));
  inv1 g276(.a(new_n290_), .O(new_n291_));
  nor2 g277(.a(new_n291_), .b(new_n289_), .O(new_n292_));
  nor2 g278(.a(new_n292_), .b(new_n284_), .O(new_n293_));
  inv1 g279(.a(new_n293_), .O(new_n294_));
  nor2 g280(.a(new_n294_), .b(new_n279_), .O(new_n295_));
  inv1 g281(.a(new_n295_), .O(new_n296_));
  nor2 g282(.a(new_n296_), .b(new_n271_), .O(new_n297_));
  inv1 g283(.a(new_n297_), .O(o_0_));
  nor2 g284(.a(new_n65_), .b(new_n24_), .O(new_n299_));
  nor2 g285(.a(new_n299_), .b(new_n51_), .O(new_n300_));
  inv1 g286(.a(new_n183_), .O(new_n301_));
  nor2 g287(.a(new_n301_), .b(new_n42_), .O(new_n302_));
  nor2 g288(.a(new_n302_), .b(new_n300_), .O(new_n303_));
  nor2 g289(.a(new_n303_), .b(i_9_), .O(new_n304_));
  nor2 g290(.a(new_n49_), .b(i_2_), .O(new_n305_));
  inv1 g291(.a(new_n305_), .O(new_n306_));
  nor2 g292(.a(new_n306_), .b(new_n53_), .O(new_n307_));
  nor2 g293(.a(new_n307_), .b(new_n234_), .O(new_n308_));
  inv1 g294(.a(new_n308_), .O(new_n309_));
  nor2 g295(.a(new_n286_), .b(new_n139_), .O(new_n310_));
  nor2 g296(.a(new_n190_), .b(new_n181_), .O(new_n311_));
  nor2 g297(.a(new_n311_), .b(new_n310_), .O(new_n312_));
  inv1 g298(.a(new_n312_), .O(new_n313_));
  nor2 g299(.a(new_n313_), .b(new_n309_), .O(new_n314_));
  inv1 g300(.a(new_n314_), .O(new_n315_));
  inv1 g301(.a(new_n267_), .O(new_n316_));
  nor2 g302(.a(new_n316_), .b(new_n252_), .O(new_n317_));
  nor2 g303(.a(new_n86_), .b(new_n22_), .O(new_n318_));
  nor2 g304(.a(new_n318_), .b(new_n317_), .O(new_n319_));
  inv1 g305(.a(new_n319_), .O(new_n320_));
  nor2 g306(.a(new_n320_), .b(new_n315_), .O(new_n321_));
  inv1 g307(.a(new_n321_), .O(new_n322_));
  nor2 g308(.a(new_n322_), .b(new_n304_), .O(new_n323_));
  inv1 g309(.a(new_n323_), .O(new_n324_));
  nor2 g310(.a(new_n324_), .b(new_n228_), .O(new_n325_));
  inv1 g311(.a(new_n325_), .O(new_n326_));
  nor2 g312(.a(new_n326_), .b(new_n220_), .O(new_n327_));
  inv1 g313(.a(new_n327_), .O(o_3_));
endmodule


