// Benchmark "top" written by ABC on Wed Jan 17 21:32:49 2024

module top ( 
    i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_,
    i_12_, i_1_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_,
    i_16_, i_22_, i_15_, i_19_,
    o_1_, o_2_, o_0_, o_7_, o_5_, o_6_, o_3_, o_4_  );
  input  i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_,
    i_4_, i_12_, i_1_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_,
    i_21_, i_16_, i_22_, i_15_, i_19_;
  output o_1_, o_2_, o_0_, o_7_, o_5_, o_6_, o_3_, o_4_;
  wire new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_;
  nor2 g000(.a(i_4_), .b(i_9_), .O(new_n34_));
  inv1 g001(.a(new_n34_), .O(new_n35_));
  nor2 g002(.a(i_11_), .b(i_12_), .O(new_n36_));
  inv1 g003(.a(new_n36_), .O(new_n37_));
  nor2 g004(.a(new_n37_), .b(new_n35_), .O(new_n38_));
  inv1 g005(.a(new_n38_), .O(new_n39_));
  nor2 g006(.a(i_16_), .b(i_14_), .O(new_n40_));
  inv1 g007(.a(new_n40_), .O(new_n41_));
  nor2 g008(.a(i_6_), .b(i_8_), .O(new_n42_));
  inv1 g009(.a(new_n42_), .O(new_n43_));
  nor2 g010(.a(i_1_), .b(i_3_), .O(new_n44_));
  inv1 g011(.a(new_n44_), .O(new_n45_));
  nor2 g012(.a(new_n45_), .b(new_n43_), .O(new_n46_));
  inv1 g013(.a(new_n46_), .O(new_n47_));
  nor2 g014(.a(new_n47_), .b(new_n41_), .O(new_n48_));
  inv1 g015(.a(new_n48_), .O(new_n49_));
  nor2 g016(.a(new_n49_), .b(new_n39_), .O(new_n50_));
  inv1 g017(.a(new_n50_), .O(new_n51_));
  nor2 g018(.a(i_22_), .b(i_23_), .O(new_n52_));
  inv1 g019(.a(new_n52_), .O(new_n53_));
  nor2 g020(.a(new_n53_), .b(i_17_), .O(new_n54_));
  inv1 g021(.a(new_n54_), .O(new_n55_));
  nor2 g022(.a(new_n55_), .b(i_20_), .O(new_n56_));
  inv1 g023(.a(new_n56_), .O(new_n57_));
  inv1 g024(.a(i_19_), .O(new_n58_));
  nor2 g025(.a(i_13_), .b(i_5_), .O(new_n59_));
  inv1 g026(.a(new_n59_), .O(new_n60_));
  nor2 g027(.a(new_n60_), .b(new_n58_), .O(new_n61_));
  inv1 g028(.a(i_24_), .O(new_n62_));
  inv1 g029(.a(i_7_), .O(new_n63_));
  inv1 g030(.a(i_13_), .O(new_n64_));
  nor2 g031(.a(new_n64_), .b(new_n63_), .O(new_n65_));
  inv1 g032(.a(new_n65_), .O(new_n66_));
  nor2 g033(.a(new_n66_), .b(new_n62_), .O(new_n67_));
  nor2 g034(.a(new_n67_), .b(new_n61_), .O(new_n68_));
  nor2 g035(.a(new_n68_), .b(new_n57_), .O(new_n69_));
  inv1 g036(.a(new_n69_), .O(new_n70_));
  nor2 g037(.a(new_n70_), .b(new_n51_), .O(new_n71_));
  nor2 g038(.a(i_24_), .b(i_10_), .O(new_n72_));
  inv1 g039(.a(new_n72_), .O(new_n73_));
  inv1 g040(.a(i_0_), .O(new_n74_));
  nor2 g041(.a(new_n74_), .b(i_2_), .O(new_n75_));
  inv1 g042(.a(new_n75_), .O(new_n76_));
  nor2 g043(.a(new_n76_), .b(new_n73_), .O(new_n77_));
  inv1 g044(.a(new_n77_), .O(new_n78_));
  nor2 g045(.a(new_n78_), .b(new_n57_), .O(new_n79_));
  inv1 g046(.a(new_n79_), .O(new_n80_));
  nor2 g047(.a(new_n80_), .b(new_n51_), .O(new_n81_));
  inv1 g048(.a(i_17_), .O(new_n82_));
  inv1 g049(.a(i_16_), .O(new_n83_));
  nor2 g050(.a(new_n83_), .b(new_n82_), .O(new_n84_));
  inv1 g051(.a(new_n84_), .O(new_n85_));
  inv1 g052(.a(i_20_), .O(new_n86_));
  inv1 g053(.a(i_14_), .O(new_n87_));
  nor2 g054(.a(new_n87_), .b(new_n86_), .O(new_n88_));
  inv1 g055(.a(new_n88_), .O(new_n89_));
  nor2 g056(.a(new_n89_), .b(new_n85_), .O(new_n90_));
  inv1 g057(.a(new_n90_), .O(new_n91_));
  inv1 g058(.a(i_3_), .O(new_n92_));
  inv1 g059(.a(i_1_), .O(new_n93_));
  nor2 g060(.a(new_n93_), .b(new_n92_), .O(new_n94_));
  inv1 g061(.a(new_n94_), .O(new_n95_));
  inv1 g062(.a(i_21_), .O(new_n96_));
  nor2 g063(.a(new_n96_), .b(i_2_), .O(new_n97_));
  inv1 g064(.a(new_n97_), .O(new_n98_));
  nor2 g065(.a(new_n98_), .b(new_n95_), .O(new_n99_));
  inv1 g066(.a(new_n99_), .O(new_n100_));
  nor2 g067(.a(new_n100_), .b(new_n91_), .O(new_n101_));
  inv1 g068(.a(new_n101_), .O(new_n102_));
  inv1 g069(.a(i_23_), .O(new_n103_));
  inv1 g070(.a(i_22_), .O(new_n104_));
  nor2 g071(.a(new_n104_), .b(new_n103_), .O(new_n105_));
  inv1 g072(.a(new_n105_), .O(new_n106_));
  nor2 g073(.a(new_n106_), .b(i_24_), .O(new_n107_));
  inv1 g074(.a(new_n107_), .O(new_n108_));
  inv1 g075(.a(i_8_), .O(new_n109_));
  inv1 g076(.a(i_6_), .O(new_n110_));
  nor2 g077(.a(new_n110_), .b(new_n109_), .O(new_n111_));
  inv1 g078(.a(new_n111_), .O(new_n112_));
  inv1 g079(.a(i_9_), .O(new_n113_));
  inv1 g080(.a(i_12_), .O(new_n114_));
  nor2 g081(.a(new_n114_), .b(new_n113_), .O(new_n115_));
  inv1 g082(.a(new_n115_), .O(new_n116_));
  nor2 g083(.a(new_n116_), .b(new_n112_), .O(new_n117_));
  inv1 g084(.a(new_n117_), .O(new_n118_));
  inv1 g085(.a(i_11_), .O(new_n119_));
  inv1 g086(.a(i_4_), .O(new_n120_));
  nor2 g087(.a(new_n120_), .b(i_10_), .O(new_n121_));
  inv1 g088(.a(new_n121_), .O(new_n122_));
  nor2 g089(.a(new_n122_), .b(new_n119_), .O(new_n123_));
  inv1 g090(.a(new_n123_), .O(new_n124_));
  nor2 g091(.a(new_n124_), .b(new_n118_), .O(new_n125_));
  inv1 g092(.a(new_n125_), .O(new_n126_));
  nor2 g093(.a(new_n126_), .b(new_n108_), .O(new_n127_));
  inv1 g094(.a(new_n127_), .O(new_n128_));
  nor2 g095(.a(new_n128_), .b(new_n102_), .O(new_n129_));
  nor2 g096(.a(new_n129_), .b(new_n81_), .O(new_n130_));
  inv1 g097(.a(new_n130_), .O(new_n131_));
  nor2 g098(.a(new_n131_), .b(new_n71_), .O(new_n132_));
  inv1 g099(.a(new_n132_), .O(new_n133_));
  inv1 g100(.a(i_18_), .O(new_n134_));
  nor2 g101(.a(new_n62_), .b(new_n134_), .O(new_n135_));
  inv1 g102(.a(new_n135_), .O(new_n136_));
  nor2 g103(.a(new_n136_), .b(new_n106_), .O(new_n137_));
  inv1 g104(.a(new_n137_), .O(new_n138_));
  nor2 g105(.a(new_n138_), .b(new_n91_), .O(new_n139_));
  inv1 g106(.a(i_15_), .O(new_n140_));
  nor2 g107(.a(new_n140_), .b(new_n64_), .O(new_n141_));
  inv1 g108(.a(new_n141_), .O(new_n142_));
  nor2 g109(.a(new_n142_), .b(new_n85_), .O(new_n143_));
  inv1 g110(.a(new_n143_), .O(new_n144_));
  nor2 g111(.a(new_n144_), .b(new_n89_), .O(new_n145_));
  inv1 g112(.a(new_n145_), .O(new_n146_));
  nor2 g113(.a(new_n146_), .b(new_n108_), .O(new_n147_));
  nor2 g114(.a(new_n147_), .b(new_n139_), .O(new_n148_));
  nor2 g115(.a(new_n112_), .b(new_n119_), .O(new_n149_));
  inv1 g116(.a(new_n149_), .O(new_n150_));
  nor2 g117(.a(new_n95_), .b(new_n120_), .O(new_n151_));
  inv1 g118(.a(new_n151_), .O(new_n152_));
  inv1 g119(.a(i_5_), .O(new_n153_));
  nor2 g120(.a(new_n116_), .b(new_n153_), .O(new_n154_));
  inv1 g121(.a(new_n154_), .O(new_n155_));
  nor2 g122(.a(new_n155_), .b(new_n152_), .O(new_n156_));
  inv1 g123(.a(new_n156_), .O(new_n157_));
  nor2 g124(.a(new_n157_), .b(new_n150_), .O(new_n158_));
  inv1 g125(.a(new_n158_), .O(new_n159_));
  nor2 g126(.a(new_n159_), .b(new_n148_), .O(new_n160_));
  nor2 g127(.a(new_n106_), .b(new_n86_), .O(new_n161_));
  inv1 g128(.a(new_n161_), .O(new_n162_));
  nor2 g129(.a(new_n119_), .b(new_n87_), .O(new_n163_));
  inv1 g130(.a(new_n163_), .O(new_n164_));
  nor2 g131(.a(new_n164_), .b(new_n85_), .O(new_n165_));
  inv1 g132(.a(new_n165_), .O(new_n166_));
  nor2 g133(.a(new_n166_), .b(new_n162_), .O(new_n167_));
  inv1 g134(.a(new_n167_), .O(new_n168_));
  nor2 g135(.a(new_n60_), .b(new_n140_), .O(new_n169_));
  inv1 g136(.a(new_n169_), .O(new_n170_));
  nor2 g137(.a(new_n170_), .b(new_n118_), .O(new_n171_));
  inv1 g138(.a(new_n171_), .O(new_n172_));
  nor2 g139(.a(new_n172_), .b(new_n168_), .O(new_n173_));
  inv1 g140(.a(new_n139_), .O(new_n174_));
  nor2 g141(.a(new_n116_), .b(new_n64_), .O(new_n175_));
  inv1 g142(.a(new_n175_), .O(new_n176_));
  nor2 g143(.a(new_n176_), .b(new_n150_), .O(new_n177_));
  inv1 g144(.a(new_n177_), .O(new_n178_));
  nor2 g145(.a(new_n178_), .b(new_n174_), .O(new_n179_));
  nor2 g146(.a(new_n179_), .b(new_n173_), .O(new_n180_));
  nor2 g147(.a(new_n180_), .b(new_n152_), .O(new_n181_));
  nor2 g148(.a(new_n64_), .b(new_n153_), .O(new_n182_));
  inv1 g149(.a(new_n182_), .O(new_n183_));
  nor2 g150(.a(new_n183_), .b(i_24_), .O(new_n184_));
  inv1 g151(.a(new_n184_), .O(new_n185_));
  nor2 g152(.a(new_n185_), .b(new_n58_), .O(new_n186_));
  inv1 g153(.a(new_n186_), .O(new_n187_));
  nor2 g154(.a(new_n187_), .b(new_n57_), .O(new_n188_));
  inv1 g155(.a(new_n188_), .O(new_n189_));
  nor2 g156(.a(new_n189_), .b(new_n51_), .O(new_n190_));
  nor2 g157(.a(new_n63_), .b(i_20_), .O(new_n191_));
  inv1 g158(.a(new_n191_), .O(new_n192_));
  nor2 g159(.a(new_n192_), .b(new_n43_), .O(new_n193_));
  inv1 g160(.a(new_n193_), .O(new_n194_));
  nor2 g161(.a(new_n194_), .b(new_n41_), .O(new_n195_));
  inv1 g162(.a(new_n195_), .O(new_n196_));
  nor2 g163(.a(i_3_), .b(new_n153_), .O(new_n197_));
  inv1 g164(.a(new_n197_), .O(new_n198_));
  nor2 g165(.a(new_n62_), .b(i_1_), .O(new_n199_));
  inv1 g166(.a(new_n199_), .O(new_n200_));
  nor2 g167(.a(new_n200_), .b(new_n198_), .O(new_n201_));
  inv1 g168(.a(new_n201_), .O(new_n202_));
  nor2 g169(.a(new_n202_), .b(new_n55_), .O(new_n203_));
  inv1 g170(.a(new_n203_), .O(new_n204_));
  nor2 g171(.a(new_n204_), .b(new_n39_), .O(new_n205_));
  inv1 g172(.a(new_n205_), .O(new_n206_));
  nor2 g173(.a(new_n206_), .b(new_n196_), .O(new_n207_));
  nor2 g174(.a(new_n207_), .b(new_n190_), .O(new_n208_));
  inv1 g175(.a(new_n208_), .O(new_n209_));
  nor2 g176(.a(new_n209_), .b(new_n181_), .O(new_n210_));
  inv1 g177(.a(new_n210_), .O(new_n211_));
  nor2 g178(.a(new_n211_), .b(new_n160_), .O(new_n212_));
  inv1 g179(.a(new_n212_), .O(new_n213_));
  nor2 g180(.a(new_n213_), .b(new_n133_), .O(new_n214_));
  inv1 g181(.a(new_n214_), .O(o_1_));
  nor2 g182(.a(new_n136_), .b(new_n64_), .O(new_n216_));
  nor2 g183(.a(new_n216_), .b(new_n169_), .O(new_n217_));
  inv1 g184(.a(new_n217_), .O(new_n218_));
  nor2 g185(.a(new_n98_), .b(new_n73_), .O(new_n219_));
  nor2 g186(.a(new_n136_), .b(new_n153_), .O(new_n220_));
  nor2 g187(.a(new_n220_), .b(new_n219_), .O(new_n221_));
  inv1 g188(.a(new_n221_), .O(new_n222_));
  nor2 g189(.a(new_n222_), .b(new_n218_), .O(new_n223_));
  inv1 g190(.a(new_n223_), .O(new_n224_));
  nor2 g191(.a(new_n185_), .b(new_n140_), .O(new_n225_));
  nor2 g192(.a(new_n225_), .b(new_n224_), .O(new_n226_));
  nor2 g193(.a(new_n110_), .b(new_n86_), .O(new_n227_));
  inv1 g194(.a(new_n227_), .O(new_n228_));
  nor2 g195(.a(new_n228_), .b(new_n95_), .O(new_n229_));
  inv1 g196(.a(new_n229_), .O(new_n230_));
  nor2 g197(.a(new_n230_), .b(new_n164_), .O(new_n231_));
  inv1 g198(.a(new_n231_), .O(new_n232_));
  nor2 g199(.a(new_n232_), .b(new_n226_), .O(o_2_));
  nor2 g200(.a(new_n186_), .b(new_n77_), .O(new_n234_));
  inv1 g201(.a(new_n234_), .O(new_n235_));
  nor2 g202(.a(new_n153_), .b(new_n63_), .O(new_n236_));
  inv1 g203(.a(new_n236_), .O(new_n237_));
  nor2 g204(.a(new_n237_), .b(new_n62_), .O(new_n238_));
  nor2 g205(.a(new_n238_), .b(new_n61_), .O(new_n239_));
  inv1 g206(.a(new_n239_), .O(new_n240_));
  nor2 g207(.a(new_n240_), .b(new_n67_), .O(new_n241_));
  inv1 g208(.a(new_n241_), .O(new_n242_));
  nor2 g209(.a(new_n242_), .b(new_n235_), .O(new_n243_));
  nor2 g210(.a(i_6_), .b(i_20_), .O(new_n244_));
  inv1 g211(.a(new_n244_), .O(new_n245_));
  nor2 g212(.a(i_3_), .b(i_14_), .O(new_n246_));
  inv1 g213(.a(new_n246_), .O(new_n247_));
  nor2 g214(.a(i_11_), .b(i_1_), .O(new_n248_));
  inv1 g215(.a(new_n248_), .O(new_n249_));
  nor2 g216(.a(new_n249_), .b(new_n247_), .O(new_n250_));
  inv1 g217(.a(new_n250_), .O(new_n251_));
  nor2 g218(.a(new_n251_), .b(new_n245_), .O(new_n252_));
  inv1 g219(.a(new_n252_), .O(new_n253_));
  nor2 g220(.a(new_n253_), .b(new_n243_), .O(o_0_));
  inv1 g221(.a(new_n226_), .O(o_7_));
  inv1 g222(.a(new_n243_), .O(o_5_));
  inv1 g223(.a(new_n219_), .O(new_n257_));
  nor2 g224(.a(new_n257_), .b(i_3_), .O(new_n258_));
  nor2 g225(.a(i_11_), .b(new_n110_), .O(new_n259_));
  inv1 g226(.a(new_n259_), .O(new_n260_));
  nor2 g227(.a(new_n260_), .b(new_n78_), .O(new_n261_));
  inv1 g228(.a(new_n67_), .O(new_n262_));
  nor2 g229(.a(i_14_), .b(new_n86_), .O(new_n263_));
  inv1 g230(.a(new_n263_), .O(new_n264_));
  nor2 g231(.a(new_n264_), .b(i_11_), .O(new_n265_));
  inv1 g232(.a(new_n265_), .O(new_n266_));
  nor2 g233(.a(new_n266_), .b(new_n262_), .O(new_n267_));
  nor2 g234(.a(new_n267_), .b(new_n261_), .O(new_n268_));
  inv1 g235(.a(new_n268_), .O(new_n269_));
  nor2 g236(.a(new_n269_), .b(new_n258_), .O(new_n270_));
  inv1 g237(.a(new_n270_), .O(new_n271_));
  nor2 g238(.a(new_n164_), .b(new_n88_), .O(new_n272_));
  nor2 g239(.a(new_n119_), .b(i_6_), .O(new_n273_));
  nor2 g240(.a(new_n273_), .b(new_n272_), .O(new_n274_));
  nor2 g241(.a(new_n274_), .b(new_n257_), .O(new_n275_));
  nor2 g242(.a(new_n273_), .b(new_n92_), .O(new_n276_));
  nor2 g243(.a(new_n276_), .b(new_n217_), .O(new_n277_));
  nor2 g244(.a(new_n277_), .b(new_n275_), .O(new_n278_));
  inv1 g245(.a(new_n278_), .O(new_n279_));
  nor2 g246(.a(new_n279_), .b(new_n271_), .O(new_n280_));
  inv1 g247(.a(new_n280_), .O(new_n281_));
  inv1 g248(.a(new_n273_), .O(new_n282_));
  nor2 g249(.a(new_n225_), .b(new_n220_), .O(new_n283_));
  nor2 g250(.a(new_n283_), .b(new_n282_), .O(new_n284_));
  nor2 g251(.a(new_n272_), .b(new_n92_), .O(new_n285_));
  nor2 g252(.a(new_n285_), .b(new_n283_), .O(new_n286_));
  nor2 g253(.a(new_n286_), .b(new_n284_), .O(new_n287_));
  inv1 g254(.a(new_n287_), .O(new_n288_));
  nor2 g255(.a(new_n288_), .b(new_n281_), .O(new_n289_));
  inv1 g256(.a(new_n289_), .O(new_n290_));
  nor2 g257(.a(new_n259_), .b(i_3_), .O(new_n291_));
  inv1 g258(.a(new_n68_), .O(new_n292_));
  nor2 g259(.a(new_n186_), .b(new_n292_), .O(new_n293_));
  inv1 g260(.a(new_n293_), .O(new_n294_));
  nor2 g261(.a(new_n294_), .b(new_n238_), .O(new_n295_));
  nor2 g262(.a(new_n295_), .b(new_n291_), .O(new_n296_));
  nor2 g263(.a(new_n266_), .b(new_n239_), .O(new_n297_));
  inv1 g264(.a(new_n272_), .O(new_n298_));
  nor2 g265(.a(new_n298_), .b(new_n217_), .O(new_n299_));
  nor2 g266(.a(new_n299_), .b(new_n297_), .O(new_n300_));
  inv1 g267(.a(new_n300_), .O(new_n301_));
  nor2 g268(.a(new_n266_), .b(new_n187_), .O(new_n302_));
  nor2 g269(.a(new_n265_), .b(i_3_), .O(new_n303_));
  nor2 g270(.a(new_n303_), .b(new_n78_), .O(new_n304_));
  nor2 g271(.a(new_n304_), .b(new_n302_), .O(new_n305_));
  inv1 g272(.a(new_n305_), .O(new_n306_));
  nor2 g273(.a(new_n306_), .b(new_n301_), .O(new_n307_));
  inv1 g274(.a(new_n307_), .O(new_n308_));
  nor2 g275(.a(new_n308_), .b(new_n296_), .O(new_n309_));
  inv1 g276(.a(new_n309_), .O(new_n310_));
  nor2 g277(.a(new_n310_), .b(new_n290_), .O(new_n311_));
  inv1 g278(.a(new_n311_), .O(o_6_));
  inv1 g279(.a(o_0_), .O(new_n313_));
  nor2 g280(.a(new_n313_), .b(i_8_), .O(new_n314_));
  nor2 g281(.a(new_n219_), .b(new_n216_), .O(new_n315_));
  nor2 g282(.a(new_n232_), .b(new_n109_), .O(new_n316_));
  inv1 g283(.a(new_n316_), .O(new_n317_));
  nor2 g284(.a(new_n317_), .b(new_n315_), .O(new_n318_));
  inv1 g285(.a(new_n283_), .O(new_n319_));
  nor2 g286(.a(new_n319_), .b(new_n169_), .O(new_n320_));
  nor2 g287(.a(new_n320_), .b(new_n317_), .O(new_n321_));
  nor2 g288(.a(new_n321_), .b(new_n318_), .O(new_n322_));
  inv1 g289(.a(new_n322_), .O(new_n323_));
  nor2 g290(.a(new_n323_), .b(new_n314_), .O(new_n324_));
  inv1 g291(.a(new_n324_), .O(o_3_));
  nor2 g292(.a(i_16_), .b(new_n120_), .O(new_n326_));
  inv1 g293(.a(new_n326_), .O(new_n327_));
  nor2 g294(.a(new_n327_), .b(new_n53_), .O(new_n328_));
  inv1 g295(.a(new_n328_), .O(new_n329_));
  nor2 g296(.a(new_n329_), .b(new_n234_), .O(new_n330_));
  nor2 g297(.a(i_16_), .b(new_n82_), .O(new_n331_));
  inv1 g298(.a(new_n331_), .O(new_n332_));
  nor2 g299(.a(new_n332_), .b(i_22_), .O(new_n333_));
  inv1 g300(.a(new_n333_), .O(new_n334_));
  nor2 g301(.a(new_n186_), .b(new_n61_), .O(new_n335_));
  nor2 g302(.a(new_n335_), .b(new_n334_), .O(new_n336_));
  nor2 g303(.a(new_n336_), .b(new_n330_), .O(new_n337_));
  inv1 g304(.a(new_n337_), .O(new_n338_));
  nor2 g305(.a(new_n225_), .b(new_n219_), .O(new_n339_));
  nor2 g306(.a(new_n339_), .b(i_8_), .O(new_n340_));
  nor2 g307(.a(new_n329_), .b(new_n241_), .O(new_n341_));
  nor2 g308(.a(new_n341_), .b(new_n340_), .O(new_n342_));
  inv1 g309(.a(new_n342_), .O(new_n343_));
  nor2 g310(.a(new_n343_), .b(new_n338_), .O(new_n344_));
  inv1 g311(.a(new_n344_), .O(new_n345_));
  nor2 g312(.a(new_n83_), .b(i_9_), .O(new_n346_));
  nor2 g313(.a(new_n83_), .b(i_4_), .O(new_n347_));
  inv1 g314(.a(new_n347_), .O(new_n348_));
  nor2 g315(.a(new_n348_), .b(new_n106_), .O(new_n349_));
  nor2 g316(.a(new_n349_), .b(new_n346_), .O(new_n350_));
  inv1 g317(.a(new_n350_), .O(new_n351_));
  nor2 g318(.a(new_n351_), .b(new_n109_), .O(new_n352_));
  nor2 g319(.a(new_n352_), .b(new_n217_), .O(new_n353_));
  nor2 g320(.a(new_n83_), .b(i_17_), .O(new_n354_));
  inv1 g321(.a(new_n354_), .O(new_n355_));
  nor2 g322(.a(new_n355_), .b(new_n104_), .O(new_n356_));
  inv1 g323(.a(new_n356_), .O(new_n357_));
  nor2 g324(.a(new_n357_), .b(new_n223_), .O(new_n358_));
  nor2 g325(.a(new_n358_), .b(new_n353_), .O(new_n359_));
  inv1 g326(.a(new_n359_), .O(new_n360_));
  nor2 g327(.a(i_16_), .b(new_n113_), .O(new_n361_));
  inv1 g328(.a(new_n361_), .O(new_n362_));
  nor2 g329(.a(new_n362_), .b(new_n293_), .O(new_n363_));
  nor2 g330(.a(new_n234_), .b(new_n109_), .O(new_n364_));
  nor2 g331(.a(new_n364_), .b(new_n363_), .O(new_n365_));
  inv1 g332(.a(new_n365_), .O(new_n366_));
  nor2 g333(.a(new_n366_), .b(new_n360_), .O(new_n367_));
  inv1 g334(.a(new_n367_), .O(new_n368_));
  inv1 g335(.a(new_n349_), .O(new_n369_));
  nor2 g336(.a(new_n369_), .b(new_n221_), .O(new_n370_));
  nor2 g337(.a(new_n334_), .b(new_n262_), .O(new_n371_));
  inv1 g338(.a(new_n346_), .O(new_n372_));
  nor2 g339(.a(new_n372_), .b(new_n257_), .O(new_n373_));
  nor2 g340(.a(new_n373_), .b(new_n371_), .O(new_n374_));
  inv1 g341(.a(new_n374_), .O(new_n375_));
  nor2 g342(.a(new_n375_), .b(new_n370_), .O(new_n376_));
  inv1 g343(.a(new_n376_), .O(new_n377_));
  nor2 g344(.a(new_n238_), .b(new_n67_), .O(new_n378_));
  nor2 g345(.a(new_n378_), .b(new_n109_), .O(new_n379_));
  nor2 g346(.a(new_n361_), .b(new_n333_), .O(new_n380_));
  nor2 g347(.a(new_n238_), .b(new_n77_), .O(new_n381_));
  nor2 g348(.a(new_n381_), .b(new_n380_), .O(new_n382_));
  nor2 g349(.a(new_n382_), .b(new_n379_), .O(new_n383_));
  inv1 g350(.a(new_n383_), .O(new_n384_));
  nor2 g351(.a(new_n384_), .b(new_n377_), .O(new_n385_));
  inv1 g352(.a(new_n385_), .O(new_n386_));
  inv1 g353(.a(new_n225_), .O(new_n387_));
  nor2 g354(.a(new_n356_), .b(new_n351_), .O(new_n388_));
  nor2 g355(.a(new_n388_), .b(new_n387_), .O(new_n389_));
  inv1 g356(.a(new_n220_), .O(new_n390_));
  nor2 g357(.a(new_n372_), .b(new_n390_), .O(new_n391_));
  inv1 g358(.a(new_n61_), .O(new_n392_));
  nor2 g359(.a(new_n392_), .b(new_n109_), .O(new_n393_));
  nor2 g360(.a(new_n390_), .b(i_8_), .O(new_n394_));
  nor2 g361(.a(new_n394_), .b(new_n393_), .O(new_n395_));
  inv1 g362(.a(new_n395_), .O(new_n396_));
  nor2 g363(.a(new_n396_), .b(new_n391_), .O(new_n397_));
  inv1 g364(.a(new_n397_), .O(new_n398_));
  nor2 g365(.a(new_n398_), .b(new_n389_), .O(new_n399_));
  inv1 g366(.a(new_n399_), .O(new_n400_));
  nor2 g367(.a(new_n400_), .b(new_n386_), .O(new_n401_));
  inv1 g368(.a(new_n401_), .O(new_n402_));
  nor2 g369(.a(new_n402_), .b(new_n368_), .O(new_n403_));
  inv1 g370(.a(new_n403_), .O(new_n404_));
  nor2 g371(.a(new_n404_), .b(new_n345_), .O(new_n405_));
  inv1 g372(.a(new_n405_), .O(o_4_));
endmodule


