// Benchmark "top" written by ABC on Wed Jan 17 21:32:50 2024

module top ( 
    i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_,
    i_12_, i_1_, i_11_, i_2_, i_18_, i_17_, i_0_, i_21_, i_16_, i_15_,
    i_19_,
    o_1_, o_19_, o_2_, o_0_, o_25_, o_12_, o_26_, o_11_, o_27_, o_14_,
    o_28_, o_13_, o_21_, o_16_, o_22_, o_15_, o_23_, o_18_, o_24_, o_17_,
    o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_  );
  input  i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_,
    i_4_, i_12_, i_1_, i_11_, i_2_, i_18_, i_17_, i_0_, i_21_, i_16_,
    i_15_, i_19_;
  output o_1_, o_19_, o_2_, o_0_, o_25_, o_12_, o_26_, o_11_, o_27_, o_14_,
    o_28_, o_13_, o_21_, o_16_, o_22_, o_15_, o_23_, o_18_, o_24_, o_17_,
    o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;
  wire new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n394_, new_n396_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n452_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_;
  inv1 g000(.a(i_18_), .O(new_n52_));
  inv1 g001(.a(i_21_), .O(new_n53_));
  nor2 g002(.a(new_n53_), .b(new_n52_), .O(new_n54_));
  inv1 g003(.a(new_n54_), .O(new_n55_));
  nor2 g004(.a(i_15_), .b(i_17_), .O(new_n56_));
  inv1 g005(.a(new_n56_), .O(new_n57_));
  nor2 g006(.a(new_n57_), .b(i_14_), .O(new_n58_));
  inv1 g007(.a(new_n58_), .O(new_n59_));
  nor2 g008(.a(new_n59_), .b(new_n55_), .O(new_n60_));
  inv1 g009(.a(new_n60_), .O(new_n61_));
  inv1 g010(.a(i_6_), .O(new_n62_));
  nor2 g011(.a(new_n62_), .b(i_5_), .O(new_n63_));
  inv1 g012(.a(new_n63_), .O(new_n64_));
  nor2 g013(.a(new_n64_), .b(i_2_), .O(new_n65_));
  inv1 g014(.a(new_n65_), .O(new_n66_));
  inv1 g015(.a(i_11_), .O(new_n67_));
  nor2 g016(.a(i_7_), .b(i_9_), .O(new_n68_));
  inv1 g017(.a(new_n68_), .O(new_n69_));
  nor2 g018(.a(new_n69_), .b(i_8_), .O(new_n70_));
  inv1 g019(.a(new_n70_), .O(new_n71_));
  nor2 g020(.a(new_n71_), .b(new_n67_), .O(new_n72_));
  inv1 g021(.a(new_n72_), .O(new_n73_));
  nor2 g022(.a(new_n73_), .b(new_n66_), .O(new_n74_));
  inv1 g023(.a(new_n74_), .O(new_n75_));
  nor2 g024(.a(new_n75_), .b(new_n61_), .O(new_n76_));
  inv1 g025(.a(i_8_), .O(new_n77_));
  nor2 g026(.a(i_5_), .b(new_n77_), .O(new_n78_));
  inv1 g027(.a(new_n78_), .O(new_n79_));
  inv1 g028(.a(i_2_), .O(new_n80_));
  nor2 g029(.a(new_n80_), .b(i_7_), .O(new_n81_));
  nor2 g030(.a(new_n81_), .b(new_n79_), .O(new_n82_));
  inv1 g031(.a(new_n82_), .O(new_n83_));
  nor2 g032(.a(new_n77_), .b(i_7_), .O(new_n84_));
  inv1 g033(.a(new_n84_), .O(new_n85_));
  nor2 g034(.a(new_n85_), .b(i_9_), .O(new_n86_));
  inv1 g035(.a(new_n86_), .O(new_n87_));
  nor2 g036(.a(new_n87_), .b(new_n83_), .O(new_n88_));
  inv1 g037(.a(new_n88_), .O(new_n89_));
  inv1 g038(.a(i_15_), .O(new_n90_));
  nor2 g039(.a(i_17_), .b(new_n52_), .O(new_n91_));
  inv1 g040(.a(new_n91_), .O(new_n92_));
  nor2 g041(.a(new_n92_), .b(new_n90_), .O(new_n93_));
  inv1 g042(.a(new_n93_), .O(new_n94_));
  nor2 g043(.a(i_21_), .b(new_n67_), .O(new_n95_));
  inv1 g044(.a(new_n95_), .O(new_n96_));
  nor2 g045(.a(new_n96_), .b(new_n94_), .O(new_n97_));
  inv1 g046(.a(new_n97_), .O(new_n98_));
  nor2 g047(.a(new_n98_), .b(new_n89_), .O(new_n99_));
  nor2 g048(.a(i_21_), .b(new_n52_), .O(new_n100_));
  inv1 g049(.a(new_n100_), .O(new_n101_));
  nor2 g050(.a(new_n101_), .b(i_17_), .O(new_n102_));
  inv1 g051(.a(new_n102_), .O(new_n103_));
  nor2 g052(.a(new_n77_), .b(i_9_), .O(new_n104_));
  inv1 g053(.a(new_n104_), .O(new_n105_));
  nor2 g054(.a(new_n105_), .b(i_4_), .O(new_n106_));
  inv1 g055(.a(new_n106_), .O(new_n107_));
  inv1 g056(.a(i_5_), .O(new_n108_));
  nor2 g057(.a(new_n108_), .b(i_7_), .O(new_n109_));
  inv1 g058(.a(new_n109_), .O(new_n110_));
  nor2 g059(.a(new_n90_), .b(i_11_), .O(new_n111_));
  inv1 g060(.a(new_n111_), .O(new_n112_));
  nor2 g061(.a(new_n112_), .b(new_n110_), .O(new_n113_));
  inv1 g062(.a(new_n113_), .O(new_n114_));
  nor2 g063(.a(new_n114_), .b(new_n107_), .O(new_n115_));
  inv1 g064(.a(new_n115_), .O(new_n116_));
  nor2 g065(.a(new_n116_), .b(new_n103_), .O(new_n117_));
  nor2 g066(.a(new_n117_), .b(new_n99_), .O(new_n118_));
  inv1 g067(.a(new_n118_), .O(new_n119_));
  nor2 g068(.a(new_n101_), .b(new_n57_), .O(new_n120_));
  inv1 g069(.a(new_n120_), .O(new_n121_));
  nor2 g070(.a(new_n121_), .b(new_n75_), .O(new_n122_));
  nor2 g071(.a(new_n122_), .b(new_n119_), .O(new_n123_));
  inv1 g072(.a(new_n123_), .O(new_n124_));
  nor2 g073(.a(new_n124_), .b(new_n76_), .O(new_n125_));
  inv1 g074(.a(new_n125_), .O(new_n126_));
  nor2 g075(.a(new_n64_), .b(new_n80_), .O(new_n127_));
  inv1 g076(.a(new_n127_), .O(new_n128_));
  nor2 g077(.a(new_n71_), .b(i_11_), .O(new_n129_));
  inv1 g078(.a(new_n129_), .O(new_n130_));
  nor2 g079(.a(new_n130_), .b(new_n128_), .O(new_n131_));
  inv1 g080(.a(new_n131_), .O(new_n132_));
  nor2 g081(.a(new_n132_), .b(new_n121_), .O(new_n133_));
  nor2 g082(.a(new_n132_), .b(new_n61_), .O(new_n134_));
  nor2 g083(.a(new_n134_), .b(new_n133_), .O(new_n135_));
  inv1 g084(.a(new_n135_), .O(new_n136_));
  inv1 g085(.a(i_13_), .O(new_n137_));
  nor2 g086(.a(new_n137_), .b(i_14_), .O(new_n138_));
  inv1 g087(.a(new_n138_), .O(new_n139_));
  nor2 g088(.a(new_n139_), .b(new_n121_), .O(new_n140_));
  inv1 g089(.a(new_n140_), .O(new_n141_));
  nor2 g090(.a(new_n141_), .b(i_10_), .O(new_n142_));
  inv1 g091(.a(new_n142_), .O(new_n143_));
  nor2 g092(.a(new_n89_), .b(new_n67_), .O(new_n144_));
  inv1 g093(.a(new_n144_), .O(new_n145_));
  nor2 g094(.a(new_n145_), .b(new_n143_), .O(new_n146_));
  nor2 g095(.a(new_n121_), .b(i_12_), .O(new_n147_));
  inv1 g096(.a(new_n147_), .O(new_n148_));
  inv1 g097(.a(i_10_), .O(new_n149_));
  nor2 g098(.a(new_n105_), .b(new_n149_), .O(new_n150_));
  inv1 g099(.a(new_n150_), .O(new_n151_));
  inv1 g100(.a(i_4_), .O(new_n152_));
  nor2 g101(.a(new_n152_), .b(i_7_), .O(new_n153_));
  inv1 g102(.a(new_n153_), .O(new_n154_));
  nor2 g103(.a(new_n154_), .b(i_5_), .O(new_n155_));
  inv1 g104(.a(new_n155_), .O(new_n156_));
  nor2 g105(.a(new_n156_), .b(new_n151_), .O(new_n157_));
  inv1 g106(.a(new_n157_), .O(new_n158_));
  nor2 g107(.a(new_n158_), .b(new_n148_), .O(new_n159_));
  inv1 g108(.a(new_n159_), .O(new_n160_));
  nor2 g109(.a(i_2_), .b(new_n67_), .O(new_n161_));
  inv1 g110(.a(new_n161_), .O(new_n162_));
  nor2 g111(.a(new_n162_), .b(new_n139_), .O(new_n163_));
  inv1 g112(.a(new_n163_), .O(new_n164_));
  nor2 g113(.a(new_n164_), .b(new_n160_), .O(new_n165_));
  nor2 g114(.a(new_n165_), .b(new_n146_), .O(new_n166_));
  inv1 g115(.a(new_n166_), .O(new_n167_));
  inv1 g116(.a(i_9_), .O(new_n168_));
  nor2 g117(.a(new_n90_), .b(new_n168_), .O(new_n169_));
  inv1 g118(.a(new_n169_), .O(new_n170_));
  nor2 g119(.a(new_n170_), .b(new_n92_), .O(new_n171_));
  inv1 g120(.a(new_n171_), .O(new_n172_));
  nor2 g121(.a(new_n172_), .b(new_n83_), .O(new_n173_));
  inv1 g122(.a(new_n173_), .O(new_n174_));
  nor2 g123(.a(new_n174_), .b(new_n85_), .O(new_n175_));
  inv1 g124(.a(i_7_), .O(new_n176_));
  nor2 g125(.a(i_5_), .b(new_n176_), .O(new_n177_));
  inv1 g126(.a(new_n177_), .O(new_n178_));
  nor2 g127(.a(i_17_), .b(i_18_), .O(new_n179_));
  inv1 g128(.a(new_n179_), .O(new_n180_));
  nor2 g129(.a(new_n180_), .b(new_n178_), .O(new_n181_));
  inv1 g130(.a(new_n181_), .O(new_n182_));
  nor2 g131(.a(new_n90_), .b(i_9_), .O(new_n183_));
  inv1 g132(.a(new_n183_), .O(new_n184_));
  nor2 g133(.a(new_n184_), .b(new_n80_), .O(new_n185_));
  inv1 g134(.a(new_n185_), .O(new_n186_));
  nor2 g135(.a(new_n186_), .b(new_n182_), .O(new_n187_));
  nor2 g136(.a(new_n187_), .b(new_n175_), .O(new_n188_));
  nor2 g137(.a(new_n188_), .b(new_n67_), .O(new_n189_));
  nor2 g138(.a(new_n189_), .b(new_n167_), .O(new_n190_));
  inv1 g139(.a(new_n190_), .O(new_n191_));
  nor2 g140(.a(new_n191_), .b(new_n136_), .O(new_n192_));
  inv1 g141(.a(new_n192_), .O(new_n193_));
  nor2 g142(.a(new_n193_), .b(new_n126_), .O(new_n194_));
  inv1 g143(.a(new_n194_), .O(o_1_));
  inv1 g144(.a(i_17_), .O(new_n196_));
  nor2 g145(.a(new_n196_), .b(i_18_), .O(new_n197_));
  inv1 g146(.a(new_n197_), .O(new_n198_));
  nor2 g147(.a(new_n198_), .b(i_15_), .O(new_n199_));
  inv1 g148(.a(new_n199_), .O(new_n200_));
  nor2 g149(.a(new_n69_), .b(i_5_), .O(new_n201_));
  inv1 g150(.a(new_n201_), .O(new_n202_));
  nor2 g151(.a(new_n202_), .b(new_n200_), .O(o_19_));
  nor2 g152(.a(new_n69_), .b(new_n66_), .O(new_n204_));
  nor2 g153(.a(i_6_), .b(i_7_), .O(new_n205_));
  inv1 g154(.a(new_n205_), .O(new_n206_));
  nor2 g155(.a(i_15_), .b(i_9_), .O(new_n207_));
  inv1 g156(.a(new_n207_), .O(new_n208_));
  nor2 g157(.a(new_n208_), .b(i_4_), .O(new_n209_));
  inv1 g158(.a(new_n209_), .O(new_n210_));
  nor2 g159(.a(new_n210_), .b(new_n206_), .O(new_n211_));
  nor2 g160(.a(new_n211_), .b(new_n204_), .O(new_n212_));
  nor2 g161(.a(new_n212_), .b(new_n92_), .O(new_n213_));
  nor2 g162(.a(new_n62_), .b(i_7_), .O(new_n214_));
  inv1 g163(.a(new_n214_), .O(new_n215_));
  nor2 g164(.a(new_n215_), .b(i_5_), .O(new_n216_));
  inv1 g165(.a(new_n216_), .O(new_n217_));
  nor2 g166(.a(i_11_), .b(i_9_), .O(new_n218_));
  inv1 g167(.a(new_n218_), .O(new_n219_));
  nor2 g168(.a(new_n219_), .b(new_n92_), .O(new_n220_));
  inv1 g169(.a(new_n220_), .O(new_n221_));
  nor2 g170(.a(new_n221_), .b(new_n217_), .O(new_n222_));
  inv1 g171(.a(i_1_), .O(new_n223_));
  nor2 g172(.a(i_17_), .b(new_n223_), .O(new_n224_));
  inv1 g173(.a(new_n224_), .O(new_n225_));
  nor2 g174(.a(new_n225_), .b(new_n178_), .O(new_n226_));
  inv1 g175(.a(new_n226_), .O(new_n227_));
  inv1 g176(.a(i_16_), .O(new_n228_));
  nor2 g177(.a(new_n228_), .b(i_18_), .O(new_n229_));
  inv1 g178(.a(new_n229_), .O(new_n230_));
  nor2 g179(.a(new_n230_), .b(new_n208_), .O(new_n231_));
  inv1 g180(.a(new_n231_), .O(new_n232_));
  nor2 g181(.a(new_n232_), .b(new_n227_), .O(new_n233_));
  nor2 g182(.a(new_n233_), .b(new_n222_), .O(new_n234_));
  inv1 g183(.a(new_n234_), .O(new_n235_));
  nor2 g184(.a(new_n92_), .b(i_15_), .O(new_n236_));
  inv1 g185(.a(new_n236_), .O(new_n237_));
  nor2 g186(.a(new_n85_), .b(i_5_), .O(new_n238_));
  inv1 g187(.a(new_n238_), .O(new_n239_));
  nor2 g188(.a(new_n239_), .b(new_n237_), .O(new_n240_));
  nor2 g189(.a(new_n178_), .b(new_n77_), .O(new_n241_));
  inv1 g190(.a(new_n241_), .O(new_n242_));
  nor2 g191(.a(new_n242_), .b(new_n172_), .O(new_n243_));
  nor2 g192(.a(new_n243_), .b(new_n240_), .O(new_n244_));
  inv1 g193(.a(new_n244_), .O(new_n245_));
  nor2 g194(.a(new_n245_), .b(new_n235_), .O(new_n246_));
  inv1 g195(.a(new_n246_), .O(new_n247_));
  nor2 g196(.a(new_n247_), .b(new_n213_), .O(new_n248_));
  inv1 g197(.a(new_n248_), .O(new_n249_));
  nor2 g198(.a(new_n85_), .b(new_n108_), .O(new_n250_));
  inv1 g199(.a(new_n250_), .O(new_n251_));
  nor2 g200(.a(new_n251_), .b(i_4_), .O(new_n252_));
  inv1 g201(.a(new_n252_), .O(new_n253_));
  inv1 g202(.a(i_12_), .O(new_n254_));
  nor2 g203(.a(new_n121_), .b(new_n254_), .O(new_n255_));
  inv1 g204(.a(new_n255_), .O(new_n256_));
  nor2 g205(.a(new_n256_), .b(new_n253_), .O(new_n257_));
  nor2 g206(.a(i_5_), .b(i_7_), .O(new_n258_));
  inv1 g207(.a(new_n258_), .O(new_n259_));
  nor2 g208(.a(new_n259_), .b(new_n80_), .O(new_n260_));
  inv1 g209(.a(new_n260_), .O(new_n261_));
  nor2 g210(.a(new_n112_), .b(new_n77_), .O(new_n262_));
  inv1 g211(.a(new_n262_), .O(new_n263_));
  nor2 g212(.a(new_n263_), .b(new_n261_), .O(new_n264_));
  inv1 g213(.a(new_n264_), .O(new_n265_));
  nor2 g214(.a(new_n265_), .b(new_n103_), .O(new_n266_));
  nor2 g215(.a(new_n266_), .b(new_n257_), .O(new_n267_));
  inv1 g216(.a(new_n267_), .O(new_n268_));
  nor2 g217(.a(i_19_), .b(new_n52_), .O(new_n269_));
  inv1 g218(.a(new_n269_), .O(new_n270_));
  nor2 g219(.a(new_n184_), .b(i_17_), .O(new_n271_));
  inv1 g220(.a(new_n271_), .O(new_n272_));
  nor2 g221(.a(new_n259_), .b(i_8_), .O(new_n273_));
  inv1 g222(.a(new_n273_), .O(new_n274_));
  nor2 g223(.a(new_n274_), .b(new_n272_), .O(new_n275_));
  inv1 g224(.a(new_n275_), .O(new_n276_));
  nor2 g225(.a(new_n276_), .b(new_n270_), .O(new_n277_));
  nor2 g226(.a(new_n272_), .b(new_n55_), .O(new_n278_));
  inv1 g227(.a(new_n278_), .O(new_n279_));
  nor2 g228(.a(new_n279_), .b(new_n251_), .O(new_n280_));
  nor2 g229(.a(new_n280_), .b(new_n277_), .O(new_n281_));
  inv1 g230(.a(new_n281_), .O(new_n282_));
  nor2 g231(.a(new_n282_), .b(new_n268_), .O(new_n283_));
  inv1 g232(.a(new_n283_), .O(new_n284_));
  nor2 g233(.a(new_n284_), .b(new_n249_), .O(new_n285_));
  inv1 g234(.a(new_n285_), .O(new_n286_));
  nor2 g235(.a(new_n265_), .b(new_n172_), .O(new_n287_));
  nor2 g236(.a(new_n254_), .b(new_n168_), .O(new_n288_));
  inv1 g237(.a(new_n288_), .O(new_n289_));
  nor2 g238(.a(new_n289_), .b(new_n237_), .O(new_n290_));
  inv1 g239(.a(new_n290_), .O(new_n291_));
  nor2 g240(.a(new_n291_), .b(new_n253_), .O(new_n292_));
  nor2 g241(.a(new_n292_), .b(new_n287_), .O(new_n293_));
  inv1 g242(.a(new_n293_), .O(new_n294_));
  nor2 g243(.a(new_n242_), .b(new_n94_), .O(new_n295_));
  inv1 g244(.a(new_n295_), .O(new_n296_));
  nor2 g245(.a(new_n296_), .b(i_9_), .O(new_n297_));
  nor2 g246(.a(new_n53_), .b(i_9_), .O(new_n298_));
  nor2 g247(.a(new_n298_), .b(new_n80_), .O(new_n299_));
  nor2 g248(.a(new_n94_), .b(new_n79_), .O(new_n300_));
  inv1 g249(.a(new_n300_), .O(new_n301_));
  nor2 g250(.a(new_n301_), .b(new_n299_), .O(new_n302_));
  nor2 g251(.a(new_n302_), .b(new_n297_), .O(new_n303_));
  inv1 g252(.a(new_n303_), .O(new_n304_));
  nor2 g253(.a(new_n304_), .b(new_n294_), .O(new_n305_));
  inv1 g254(.a(new_n305_), .O(new_n306_));
  nor2 g255(.a(new_n110_), .b(i_8_), .O(new_n307_));
  inv1 g256(.a(new_n307_), .O(new_n308_));
  nor2 g257(.a(new_n57_), .b(i_9_), .O(new_n309_));
  inv1 g258(.a(new_n309_), .O(new_n310_));
  inv1 g259(.a(i_19_), .O(new_n311_));
  nor2 g260(.a(new_n311_), .b(new_n52_), .O(new_n312_));
  inv1 g261(.a(new_n312_), .O(new_n313_));
  nor2 g262(.a(new_n313_), .b(new_n310_), .O(new_n314_));
  inv1 g263(.a(new_n314_), .O(new_n315_));
  nor2 g264(.a(new_n315_), .b(new_n308_), .O(new_n316_));
  nor2 g265(.a(new_n308_), .b(new_n270_), .O(new_n317_));
  inv1 g266(.a(new_n317_), .O(new_n318_));
  nor2 g267(.a(new_n318_), .b(new_n310_), .O(new_n319_));
  nor2 g268(.a(new_n319_), .b(new_n316_), .O(new_n320_));
  inv1 g269(.a(new_n320_), .O(new_n321_));
  nor2 g270(.a(new_n276_), .b(new_n52_), .O(new_n322_));
  inv1 g271(.a(new_n322_), .O(new_n323_));
  nor2 g272(.a(new_n323_), .b(new_n311_), .O(new_n324_));
  nor2 g273(.a(new_n324_), .b(new_n321_), .O(new_n325_));
  inv1 g274(.a(new_n325_), .O(new_n326_));
  nor2 g275(.a(i_18_), .b(i_9_), .O(new_n327_));
  inv1 g276(.a(new_n327_), .O(new_n328_));
  nor2 g277(.a(new_n328_), .b(i_15_), .O(new_n329_));
  inv1 g278(.a(new_n329_), .O(new_n330_));
  nor2 g279(.a(new_n330_), .b(new_n227_), .O(o_11_));
  inv1 g280(.a(o_11_), .O(new_n332_));
  nor2 g281(.a(new_n332_), .b(new_n77_), .O(new_n333_));
  nor2 g282(.a(new_n333_), .b(new_n117_), .O(new_n334_));
  inv1 g283(.a(new_n334_), .O(new_n335_));
  nor2 g284(.a(new_n108_), .b(new_n77_), .O(new_n336_));
  inv1 g285(.a(new_n336_), .O(new_n337_));
  nor2 g286(.a(new_n337_), .b(new_n237_), .O(new_n338_));
  inv1 g287(.a(new_n338_), .O(new_n339_));
  nor2 g288(.a(new_n254_), .b(i_7_), .O(new_n340_));
  inv1 g289(.a(new_n340_), .O(new_n341_));
  nor2 g290(.a(new_n341_), .b(new_n298_), .O(new_n342_));
  nor2 g291(.a(new_n342_), .b(new_n339_), .O(new_n343_));
  nor2 g292(.a(new_n237_), .b(new_n69_), .O(new_n344_));
  inv1 g293(.a(new_n344_), .O(new_n345_));
  nor2 g294(.a(i_12_), .b(i_6_), .O(new_n346_));
  inv1 g295(.a(new_n346_), .O(new_n347_));
  nor2 g296(.a(new_n347_), .b(new_n345_), .O(new_n348_));
  nor2 g297(.a(new_n348_), .b(new_n343_), .O(new_n349_));
  inv1 g298(.a(new_n349_), .O(new_n350_));
  nor2 g299(.a(new_n350_), .b(new_n335_), .O(new_n351_));
  inv1 g300(.a(new_n351_), .O(new_n352_));
  nor2 g301(.a(new_n352_), .b(new_n326_), .O(new_n353_));
  inv1 g302(.a(new_n353_), .O(new_n354_));
  nor2 g303(.a(new_n354_), .b(new_n306_), .O(new_n355_));
  inv1 g304(.a(new_n355_), .O(new_n356_));
  nor2 g305(.a(new_n356_), .b(new_n286_), .O(new_n357_));
  inv1 g306(.a(new_n357_), .O(o_2_));
  nor2 g307(.a(new_n176_), .b(i_9_), .O(new_n359_));
  inv1 g308(.a(new_n359_), .O(new_n360_));
  nor2 g309(.a(new_n360_), .b(i_5_), .O(new_n361_));
  inv1 g310(.a(new_n361_), .O(new_n362_));
  nor2 g311(.a(new_n198_), .b(new_n184_), .O(new_n363_));
  inv1 g312(.a(new_n363_), .O(new_n364_));
  nor2 g313(.a(new_n364_), .b(new_n362_), .O(new_n365_));
  nor2 g314(.a(new_n208_), .b(new_n108_), .O(new_n366_));
  inv1 g315(.a(new_n366_), .O(new_n367_));
  nor2 g316(.a(new_n367_), .b(new_n198_), .O(new_n368_));
  nor2 g317(.a(new_n368_), .b(o_19_), .O(new_n369_));
  inv1 g318(.a(new_n369_), .O(new_n370_));
  nor2 g319(.a(new_n370_), .b(new_n365_), .O(new_n371_));
  inv1 g320(.a(new_n371_), .O(new_n372_));
  nor2 g321(.a(new_n259_), .b(i_0_), .O(new_n373_));
  inv1 g322(.a(new_n373_), .O(new_n374_));
  nor2 g323(.a(new_n374_), .b(new_n364_), .O(new_n375_));
  nor2 g324(.a(new_n110_), .b(i_9_), .O(new_n376_));
  inv1 g325(.a(new_n376_), .O(new_n377_));
  nor2 g326(.a(new_n377_), .b(new_n198_), .O(new_n378_));
  nor2 g327(.a(new_n378_), .b(new_n375_), .O(new_n379_));
  inv1 g328(.a(new_n379_), .O(new_n380_));
  nor2 g329(.a(new_n180_), .b(i_21_), .O(new_n381_));
  inv1 g330(.a(new_n381_), .O(new_n382_));
  nor2 g331(.a(new_n254_), .b(i_14_), .O(new_n383_));
  inv1 g332(.a(new_n383_), .O(new_n384_));
  nor2 g333(.a(new_n384_), .b(new_n208_), .O(new_n385_));
  inv1 g334(.a(new_n385_), .O(new_n386_));
  nor2 g335(.a(new_n386_), .b(new_n382_), .O(new_n387_));
  inv1 g336(.a(new_n387_), .O(new_n388_));
  nor2 g337(.a(new_n388_), .b(new_n156_), .O(new_n389_));
  nor2 g338(.a(new_n389_), .b(new_n380_), .O(new_n390_));
  inv1 g339(.a(new_n390_), .O(new_n391_));
  nor2 g340(.a(new_n391_), .b(new_n372_), .O(new_n392_));
  inv1 g341(.a(new_n392_), .O(o_0_));
  inv1 g342(.a(new_n240_), .O(new_n394_));
  nor2 g343(.a(new_n394_), .b(new_n168_), .O(o_23_));
  nor2 g344(.a(o_23_), .b(new_n322_), .O(new_n396_));
  inv1 g345(.a(new_n396_), .O(o_25_));
  nor2 g346(.a(new_n362_), .b(new_n200_), .O(new_n398_));
  inv1 g347(.a(i_0_), .O(new_n399_));
  nor2 g348(.a(new_n259_), .b(new_n399_), .O(new_n400_));
  inv1 g349(.a(new_n400_), .O(new_n401_));
  nor2 g350(.a(new_n401_), .b(new_n364_), .O(new_n402_));
  nor2 g351(.a(new_n402_), .b(new_n398_), .O(new_n403_));
  inv1 g352(.a(new_n403_), .O(new_n404_));
  nor2 g353(.a(new_n404_), .b(new_n99_), .O(new_n405_));
  inv1 g354(.a(new_n405_), .O(new_n406_));
  nor2 g355(.a(i_13_), .b(i_14_), .O(new_n407_));
  inv1 g356(.a(new_n407_), .O(new_n408_));
  nor2 g357(.a(new_n408_), .b(new_n160_), .O(new_n409_));
  nor2 g358(.a(new_n409_), .b(new_n406_), .O(new_n410_));
  inv1 g359(.a(new_n410_), .O(new_n411_));
  nor2 g360(.a(new_n411_), .b(new_n167_), .O(new_n412_));
  inv1 g361(.a(new_n412_), .O(new_n413_));
  nor2 g362(.a(new_n105_), .b(new_n152_), .O(new_n414_));
  inv1 g363(.a(new_n414_), .O(new_n415_));
  nor2 g364(.a(new_n415_), .b(new_n110_), .O(new_n416_));
  inv1 g365(.a(new_n416_), .O(new_n417_));
  nor2 g366(.a(new_n417_), .b(new_n148_), .O(new_n418_));
  nor2 g367(.a(new_n418_), .b(new_n122_), .O(new_n419_));
  inv1 g368(.a(new_n419_), .O(new_n420_));
  nor2 g369(.a(i_6_), .b(i_5_), .O(new_n421_));
  inv1 g370(.a(new_n421_), .O(new_n422_));
  nor2 g371(.a(new_n422_), .b(i_4_), .O(new_n423_));
  inv1 g372(.a(new_n423_), .O(new_n424_));
  nor2 g373(.a(new_n424_), .b(new_n71_), .O(new_n425_));
  inv1 g374(.a(new_n425_), .O(new_n426_));
  nor2 g375(.a(new_n426_), .b(new_n256_), .O(new_n427_));
  nor2 g376(.a(new_n422_), .b(new_n152_), .O(new_n428_));
  inv1 g377(.a(new_n428_), .O(new_n429_));
  nor2 g378(.a(new_n429_), .b(new_n71_), .O(new_n430_));
  inv1 g379(.a(new_n430_), .O(new_n431_));
  nor2 g380(.a(new_n431_), .b(new_n148_), .O(new_n432_));
  nor2 g381(.a(new_n432_), .b(new_n427_), .O(new_n433_));
  inv1 g382(.a(new_n433_), .O(new_n434_));
  nor2 g383(.a(i_10_), .b(i_9_), .O(new_n435_));
  inv1 g384(.a(new_n435_), .O(new_n436_));
  nor2 g385(.a(new_n436_), .b(new_n408_), .O(new_n437_));
  inv1 g386(.a(new_n437_), .O(new_n438_));
  nor2 g387(.a(new_n438_), .b(new_n121_), .O(new_n439_));
  inv1 g388(.a(new_n439_), .O(new_n440_));
  nor2 g389(.a(new_n440_), .b(new_n239_), .O(new_n441_));
  nor2 g390(.a(new_n441_), .b(new_n117_), .O(new_n442_));
  inv1 g391(.a(new_n442_), .O(new_n443_));
  nor2 g392(.a(new_n443_), .b(new_n133_), .O(new_n444_));
  inv1 g393(.a(new_n444_), .O(new_n445_));
  nor2 g394(.a(new_n445_), .b(new_n434_), .O(new_n446_));
  inv1 g395(.a(new_n446_), .O(new_n447_));
  nor2 g396(.a(new_n447_), .b(new_n420_), .O(new_n448_));
  inv1 g397(.a(new_n448_), .O(new_n449_));
  nor2 g398(.a(new_n449_), .b(new_n413_), .O(new_n450_));
  inv1 g399(.a(new_n450_), .O(o_12_));
  nor2 g400(.a(i_21_), .b(i_14_), .O(new_n452_));
  nor2 g401(.a(new_n452_), .b(i_20_), .O(o_26_));
  inv1 g402(.a(i_3_), .O(new_n454_));
  inv1 g403(.a(o_23_), .O(new_n455_));
  nor2 g404(.a(new_n455_), .b(new_n454_), .O(new_n456_));
  nor2 g405(.a(new_n456_), .b(new_n297_), .O(new_n457_));
  nor2 g406(.a(new_n457_), .b(new_n311_), .O(new_n458_));
  nor2 g407(.a(new_n427_), .b(new_n316_), .O(new_n459_));
  inv1 g408(.a(new_n459_), .O(new_n460_));
  nor2 g409(.a(new_n460_), .b(new_n133_), .O(new_n461_));
  inv1 g410(.a(new_n461_), .O(new_n462_));
  nor2 g411(.a(new_n339_), .b(new_n176_), .O(new_n463_));
  inv1 g412(.a(new_n463_), .O(new_n464_));
  nor2 g413(.a(new_n464_), .b(new_n315_), .O(new_n465_));
  nor2 g414(.a(new_n404_), .b(new_n117_), .O(new_n466_));
  inv1 g415(.a(new_n466_), .O(new_n467_));
  nor2 g416(.a(new_n467_), .b(new_n465_), .O(new_n468_));
  inv1 g417(.a(new_n468_), .O(new_n469_));
  nor2 g418(.a(new_n469_), .b(new_n462_), .O(new_n470_));
  inv1 g419(.a(new_n470_), .O(new_n471_));
  nor2 g420(.a(new_n471_), .b(new_n458_), .O(new_n472_));
  inv1 g421(.a(new_n472_), .O(o_27_));
  nor2 g422(.a(i_12_), .b(new_n168_), .O(new_n474_));
  inv1 g423(.a(new_n474_), .O(new_n475_));
  nor2 g424(.a(new_n475_), .b(new_n339_), .O(new_n476_));
  inv1 g425(.a(new_n476_), .O(new_n477_));
  nor2 g426(.a(new_n477_), .b(new_n154_), .O(new_n478_));
  nor2 g427(.a(new_n418_), .b(new_n389_), .O(new_n479_));
  inv1 g428(.a(new_n479_), .O(new_n480_));
  nor2 g429(.a(new_n480_), .b(new_n406_), .O(new_n481_));
  inv1 g430(.a(new_n481_), .O(new_n482_));
  nor2 g431(.a(new_n482_), .b(new_n478_), .O(new_n483_));
  inv1 g432(.a(new_n483_), .O(new_n484_));
  nor2 g433(.a(new_n463_), .b(new_n295_), .O(new_n485_));
  nor2 g434(.a(new_n485_), .b(i_19_), .O(new_n486_));
  nor2 g435(.a(new_n375_), .b(new_n365_), .O(new_n487_));
  inv1 g436(.a(new_n487_), .O(new_n488_));
  nor2 g437(.a(new_n180_), .b(new_n112_), .O(new_n489_));
  inv1 g438(.a(new_n489_), .O(new_n490_));
  nor2 g439(.a(new_n490_), .b(new_n362_), .O(new_n491_));
  nor2 g440(.a(new_n184_), .b(i_2_), .O(new_n492_));
  inv1 g441(.a(new_n492_), .O(new_n493_));
  nor2 g442(.a(new_n493_), .b(new_n182_), .O(new_n494_));
  nor2 g443(.a(new_n494_), .b(new_n491_), .O(new_n495_));
  inv1 g444(.a(new_n495_), .O(new_n496_));
  nor2 g445(.a(new_n178_), .b(i_1_), .O(new_n497_));
  inv1 g446(.a(new_n497_), .O(new_n498_));
  nor2 g447(.a(new_n498_), .b(new_n328_), .O(new_n499_));
  nor2 g448(.a(new_n499_), .b(new_n496_), .O(new_n500_));
  inv1 g449(.a(new_n500_), .O(new_n501_));
  nor2 g450(.a(new_n501_), .b(new_n488_), .O(new_n502_));
  inv1 g451(.a(new_n502_), .O(new_n503_));
  nor2 g452(.a(new_n503_), .b(new_n189_), .O(new_n504_));
  inv1 g453(.a(new_n504_), .O(new_n505_));
  nor2 g454(.a(new_n505_), .b(new_n486_), .O(new_n506_));
  inv1 g455(.a(new_n506_), .O(new_n507_));
  nor2 g456(.a(new_n507_), .b(new_n484_), .O(new_n508_));
  inv1 g457(.a(new_n508_), .O(o_14_));
  nor2 g458(.a(new_n206_), .b(i_5_), .O(new_n510_));
  inv1 g459(.a(new_n510_), .O(new_n511_));
  nor2 g460(.a(new_n384_), .b(i_13_), .O(new_n512_));
  inv1 g461(.a(new_n512_), .O(new_n513_));
  nor2 g462(.a(new_n513_), .b(new_n151_), .O(new_n514_));
  inv1 g463(.a(new_n514_), .O(new_n515_));
  nor2 g464(.a(new_n515_), .b(new_n511_), .O(new_n516_));
  inv1 g465(.a(new_n516_), .O(new_n517_));
  nor2 g466(.a(new_n121_), .b(new_n228_), .O(new_n518_));
  inv1 g467(.a(new_n518_), .O(new_n519_));
  nor2 g468(.a(new_n519_), .b(new_n517_), .O(new_n520_));
  nor2 g469(.a(new_n121_), .b(i_16_), .O(new_n521_));
  inv1 g470(.a(new_n521_), .O(new_n522_));
  nor2 g471(.a(new_n515_), .b(new_n217_), .O(new_n523_));
  inv1 g472(.a(new_n523_), .O(new_n524_));
  nor2 g473(.a(new_n524_), .b(new_n522_), .O(new_n525_));
  nor2 g474(.a(new_n525_), .b(new_n520_), .O(new_n526_));
  inv1 g475(.a(new_n526_), .O(new_n527_));
  nor2 g476(.a(new_n61_), .b(i_12_), .O(new_n528_));
  inv1 g477(.a(new_n528_), .O(new_n529_));
  nor2 g478(.a(new_n529_), .b(new_n431_), .O(new_n530_));
  nor2 g479(.a(new_n530_), .b(new_n76_), .O(new_n531_));
  inv1 g480(.a(new_n531_), .O(new_n532_));
  nor2 g481(.a(new_n522_), .b(new_n517_), .O(new_n533_));
  nor2 g482(.a(new_n524_), .b(new_n519_), .O(new_n534_));
  nor2 g483(.a(new_n534_), .b(new_n533_), .O(new_n535_));
  inv1 g484(.a(new_n535_), .O(new_n536_));
  nor2 g485(.a(new_n536_), .b(new_n532_), .O(new_n537_));
  inv1 g486(.a(new_n537_), .O(new_n538_));
  nor2 g487(.a(new_n538_), .b(new_n527_), .O(new_n539_));
  inv1 g488(.a(new_n539_), .O(new_n540_));
  nor2 g489(.a(i_19_), .b(i_5_), .O(new_n541_));
  inv1 g490(.a(new_n541_), .O(new_n542_));
  nor2 g491(.a(new_n542_), .b(new_n364_), .O(new_n543_));
  nor2 g492(.a(new_n402_), .b(new_n243_), .O(new_n544_));
  inv1 g493(.a(new_n544_), .O(new_n545_));
  nor2 g494(.a(new_n545_), .b(new_n543_), .O(new_n546_));
  inv1 g495(.a(new_n546_), .O(new_n547_));
  nor2 g496(.a(new_n496_), .b(new_n380_), .O(new_n548_));
  inv1 g497(.a(new_n548_), .O(new_n549_));
  nor2 g498(.a(new_n549_), .b(new_n547_), .O(new_n550_));
  inv1 g499(.a(new_n550_), .O(new_n551_));
  nor2 g500(.a(new_n384_), .b(new_n67_), .O(new_n552_));
  inv1 g501(.a(new_n552_), .O(new_n553_));
  nor2 g502(.a(new_n103_), .b(new_n149_), .O(new_n554_));
  inv1 g503(.a(new_n554_), .O(new_n555_));
  nor2 g504(.a(new_n555_), .b(new_n553_), .O(new_n556_));
  inv1 g505(.a(new_n556_), .O(new_n557_));
  nor2 g506(.a(new_n557_), .b(new_n89_), .O(new_n558_));
  nor2 g507(.a(new_n558_), .b(new_n282_), .O(new_n559_));
  inv1 g508(.a(new_n559_), .O(new_n560_));
  nor2 g509(.a(new_n560_), .b(new_n551_), .O(new_n561_));
  inv1 g510(.a(new_n561_), .O(new_n562_));
  nor2 g511(.a(new_n151_), .b(new_n254_), .O(new_n563_));
  inv1 g512(.a(new_n563_), .O(new_n564_));
  nor2 g513(.a(new_n564_), .b(new_n261_), .O(new_n565_));
  inv1 g514(.a(new_n565_), .O(new_n566_));
  nor2 g515(.a(new_n566_), .b(new_n141_), .O(new_n567_));
  nor2 g516(.a(new_n567_), .b(new_n268_), .O(new_n568_));
  inv1 g517(.a(new_n568_), .O(new_n569_));
  nor2 g518(.a(new_n569_), .b(new_n306_), .O(new_n570_));
  inv1 g519(.a(new_n570_), .O(new_n571_));
  nor2 g520(.a(new_n571_), .b(new_n562_), .O(new_n572_));
  inv1 g521(.a(new_n572_), .O(new_n573_));
  nor2 g522(.a(new_n573_), .b(new_n540_), .O(new_n574_));
  inv1 g523(.a(new_n574_), .O(o_28_));
  nor2 g524(.a(new_n378_), .b(o_19_), .O(new_n576_));
  inv1 g525(.a(new_n576_), .O(new_n577_));
  nor2 g526(.a(new_n577_), .b(new_n404_), .O(new_n578_));
  inv1 g527(.a(new_n578_), .O(new_n579_));
  nor2 g528(.a(new_n579_), .b(new_n488_), .O(new_n580_));
  inv1 g529(.a(new_n580_), .O(o_13_));
  nor2 g530(.a(new_n92_), .b(i_8_), .O(new_n582_));
  inv1 g531(.a(new_n582_), .O(new_n583_));
  nor2 g532(.a(new_n583_), .b(new_n367_), .O(new_n584_));
  inv1 g533(.a(new_n584_), .O(new_n585_));
  nor2 g534(.a(new_n585_), .b(new_n215_), .O(new_n586_));
  nor2 g535(.a(o_23_), .b(new_n295_), .O(new_n587_));
  inv1 g536(.a(new_n587_), .O(new_n588_));
  nor2 g537(.a(new_n588_), .b(new_n586_), .O(new_n589_));
  nor2 g538(.a(new_n589_), .b(new_n215_), .O(new_n590_));
  nor2 g539(.a(new_n583_), .b(new_n184_), .O(new_n591_));
  inv1 g540(.a(new_n591_), .O(new_n592_));
  nor2 g541(.a(new_n592_), .b(new_n511_), .O(new_n593_));
  nor2 g542(.a(new_n593_), .b(new_n297_), .O(new_n594_));
  inv1 g543(.a(new_n594_), .O(new_n595_));
  nor2 g544(.a(new_n595_), .b(new_n590_), .O(new_n596_));
  inv1 g545(.a(new_n596_), .O(o_21_));
  nor2 g546(.a(new_n522_), .b(new_n66_), .O(new_n598_));
  nor2 g547(.a(new_n422_), .b(i_2_), .O(new_n599_));
  inv1 g548(.a(new_n599_), .O(new_n600_));
  nor2 g549(.a(new_n600_), .b(new_n519_), .O(new_n601_));
  nor2 g550(.a(new_n601_), .b(new_n598_), .O(new_n602_));
  nor2 g551(.a(new_n553_), .b(new_n87_), .O(new_n603_));
  inv1 g552(.a(new_n603_), .O(new_n604_));
  nor2 g553(.a(new_n604_), .b(new_n602_), .O(new_n605_));
  nor2 g554(.a(new_n143_), .b(new_n87_), .O(new_n606_));
  inv1 g555(.a(new_n606_), .O(new_n607_));
  nor2 g556(.a(new_n607_), .b(new_n128_), .O(new_n608_));
  nor2 g557(.a(new_n394_), .b(i_19_), .O(new_n609_));
  nor2 g558(.a(new_n609_), .b(new_n463_), .O(new_n610_));
  nor2 g559(.a(new_n610_), .b(new_n168_), .O(new_n611_));
  nor2 g560(.a(new_n611_), .b(new_n608_), .O(new_n612_));
  inv1 g561(.a(new_n612_), .O(new_n613_));
  nor2 g562(.a(new_n613_), .b(new_n605_), .O(new_n614_));
  inv1 g563(.a(new_n614_), .O(new_n615_));
  nor2 g564(.a(new_n441_), .b(new_n173_), .O(new_n616_));
  inv1 g565(.a(new_n616_), .O(new_n617_));
  nor2 g566(.a(new_n617_), .b(new_n476_), .O(new_n618_));
  inv1 g567(.a(new_n618_), .O(new_n619_));
  nor2 g568(.a(new_n152_), .b(i_14_), .O(new_n620_));
  inv1 g569(.a(new_n620_), .O(new_n621_));
  nor2 g570(.a(new_n621_), .b(new_n87_), .O(new_n622_));
  inv1 g571(.a(new_n622_), .O(new_n623_));
  nor2 g572(.a(new_n623_), .b(new_n128_), .O(new_n624_));
  inv1 g573(.a(new_n624_), .O(new_n625_));
  nor2 g574(.a(new_n625_), .b(new_n148_), .O(new_n626_));
  nor2 g575(.a(new_n626_), .b(new_n409_), .O(new_n627_));
  inv1 g576(.a(new_n627_), .O(new_n628_));
  nor2 g577(.a(new_n628_), .b(new_n619_), .O(new_n629_));
  inv1 g578(.a(new_n629_), .O(new_n630_));
  nor2 g579(.a(new_n527_), .b(new_n167_), .O(new_n631_));
  inv1 g580(.a(new_n631_), .O(new_n632_));
  nor2 g581(.a(new_n632_), .b(new_n630_), .O(new_n633_));
  inv1 g582(.a(new_n633_), .O(new_n634_));
  nor2 g583(.a(new_n634_), .b(new_n615_), .O(new_n635_));
  inv1 g584(.a(new_n635_), .O(o_16_));
  inv1 g585(.a(new_n589_), .O(new_n637_));
  nor2 g586(.a(new_n592_), .b(new_n217_), .O(new_n638_));
  nor2 g587(.a(new_n638_), .b(new_n637_), .O(new_n639_));
  inv1 g588(.a(new_n639_), .O(o_22_));
  inv1 g589(.a(new_n368_), .O(new_n641_));
  nor2 g590(.a(new_n641_), .b(i_7_), .O(o_15_));
  nor2 g591(.a(new_n422_), .b(new_n80_), .O(new_n643_));
  inv1 g592(.a(new_n643_), .O(new_n644_));
  nor2 g593(.a(new_n644_), .b(new_n607_), .O(new_n645_));
  nor2 g594(.a(new_n645_), .b(new_n536_), .O(new_n646_));
  inv1 g595(.a(new_n646_), .O(new_n647_));
  nor2 g596(.a(new_n61_), .b(new_n254_), .O(new_n648_));
  inv1 g597(.a(new_n648_), .O(new_n649_));
  nor2 g598(.a(new_n649_), .b(new_n426_), .O(new_n650_));
  nor2 g599(.a(new_n650_), .b(new_n647_), .O(new_n651_));
  inv1 g600(.a(new_n651_), .O(new_n652_));
  nor2 g601(.a(new_n324_), .b(new_n134_), .O(new_n653_));
  inv1 g602(.a(new_n653_), .O(new_n654_));
  nor2 g603(.a(new_n654_), .b(new_n652_), .O(new_n655_));
  inv1 g604(.a(new_n655_), .O(o_18_));
  nor2 g605(.a(new_n345_), .b(new_n274_), .O(new_n657_));
  nor2 g606(.a(new_n657_), .b(new_n333_), .O(new_n658_));
  inv1 g607(.a(new_n658_), .O(new_n659_));
  nor2 g608(.a(new_n659_), .b(new_n119_), .O(new_n660_));
  inv1 g609(.a(new_n660_), .O(new_n661_));
  nor2 g610(.a(new_n661_), .b(new_n480_), .O(new_n662_));
  inv1 g611(.a(new_n662_), .O(o_24_));
  nor2 g612(.a(new_n467_), .b(new_n427_), .O(new_n664_));
  inv1 g613(.a(new_n664_), .O(new_n665_));
  nor2 g614(.a(new_n665_), .b(new_n650_), .O(new_n666_));
  inv1 g615(.a(new_n666_), .O(new_n667_));
  nor2 g616(.a(new_n667_), .b(new_n136_), .O(new_n668_));
  inv1 g617(.a(new_n668_), .O(o_17_));
  nor2 g618(.a(new_n480_), .b(new_n478_), .O(new_n670_));
  inv1 g619(.a(new_n670_), .O(new_n671_));
  nor2 g620(.a(new_n650_), .b(new_n530_), .O(new_n672_));
  inv1 g621(.a(new_n672_), .O(new_n673_));
  nor2 g622(.a(new_n673_), .b(new_n671_), .O(new_n674_));
  inv1 g623(.a(new_n674_), .O(new_n675_));
  nor2 g624(.a(new_n165_), .b(new_n117_), .O(new_n676_));
  inv1 g625(.a(new_n676_), .O(new_n677_));
  nor2 g626(.a(new_n434_), .b(new_n409_), .O(new_n678_));
  inv1 g627(.a(new_n678_), .O(new_n679_));
  nor2 g628(.a(new_n679_), .b(new_n677_), .O(new_n680_));
  inv1 g629(.a(new_n680_), .O(new_n681_));
  nor2 g630(.a(new_n681_), .b(new_n675_), .O(new_n682_));
  inv1 g631(.a(new_n682_), .O(o_20_));
  nor2 g632(.a(new_n463_), .b(o_23_), .O(new_n684_));
  inv1 g633(.a(new_n684_), .O(new_n685_));
  nor2 g634(.a(new_n585_), .b(new_n206_), .O(new_n686_));
  nor2 g635(.a(new_n686_), .b(new_n593_), .O(new_n687_));
  inv1 g636(.a(new_n687_), .O(new_n688_));
  nor2 g637(.a(new_n688_), .b(new_n685_), .O(new_n689_));
  inv1 g638(.a(new_n689_), .O(new_n690_));
  nor2 g639(.a(new_n690_), .b(o_13_), .O(new_n691_));
  inv1 g640(.a(new_n691_), .O(o_10_));
  nor2 g641(.a(new_n319_), .b(o_19_), .O(new_n693_));
  inv1 g642(.a(new_n693_), .O(new_n694_));
  nor2 g643(.a(new_n343_), .b(new_n280_), .O(new_n695_));
  inv1 g644(.a(new_n695_), .O(new_n696_));
  nor2 g645(.a(new_n696_), .b(new_n694_), .O(new_n697_));
  inv1 g646(.a(new_n697_), .O(new_n698_));
  nor2 g647(.a(new_n294_), .b(new_n122_), .O(new_n699_));
  inv1 g648(.a(new_n699_), .O(new_n700_));
  nor2 g649(.a(new_n700_), .b(new_n698_), .O(new_n701_));
  inv1 g650(.a(new_n701_), .O(new_n702_));
  nor2 g651(.a(new_n432_), .b(new_n389_), .O(new_n703_));
  inv1 g652(.a(new_n703_), .O(new_n704_));
  inv1 g653(.a(new_n81_), .O(new_n705_));
  nor2 g654(.a(new_n705_), .b(i_12_), .O(new_n706_));
  inv1 g655(.a(new_n706_), .O(new_n707_));
  nor2 g656(.a(new_n707_), .b(new_n415_), .O(new_n708_));
  inv1 g657(.a(new_n708_), .O(new_n709_));
  nor2 g658(.a(new_n709_), .b(new_n141_), .O(new_n710_));
  nor2 g659(.a(new_n710_), .b(o_15_), .O(new_n711_));
  inv1 g660(.a(new_n711_), .O(new_n712_));
  nor2 g661(.a(new_n712_), .b(new_n704_), .O(new_n713_));
  inv1 g662(.a(new_n713_), .O(new_n714_));
  nor2 g663(.a(new_n714_), .b(new_n569_), .O(new_n715_));
  inv1 g664(.a(new_n715_), .O(new_n716_));
  nor2 g665(.a(new_n645_), .b(new_n608_), .O(new_n717_));
  inv1 g666(.a(new_n717_), .O(new_n718_));
  nor2 g667(.a(new_n718_), .b(new_n716_), .O(new_n719_));
  inv1 g668(.a(new_n719_), .O(new_n720_));
  nor2 g669(.a(new_n720_), .b(new_n702_), .O(new_n721_));
  inv1 g670(.a(new_n721_), .O(o_9_));
  nor2 g671(.a(new_n485_), .b(i_9_), .O(new_n723_));
  nor2 g672(.a(new_n455_), .b(new_n228_), .O(new_n724_));
  nor2 g673(.a(new_n724_), .b(new_n277_), .O(new_n725_));
  inv1 g674(.a(new_n725_), .O(new_n726_));
  nor2 g675(.a(new_n726_), .b(new_n326_), .O(new_n727_));
  inv1 g676(.a(new_n727_), .O(new_n728_));
  nor2 g677(.a(new_n728_), .b(new_n723_), .O(new_n729_));
  inv1 g678(.a(new_n729_), .O(o_7_));
  inv1 g679(.a(i_14_), .O(new_n731_));
  nor2 g680(.a(new_n731_), .b(i_20_), .O(o_8_));
  nor2 g681(.a(new_n532_), .b(new_n134_), .O(new_n733_));
  inv1 g682(.a(new_n733_), .O(new_n734_));
  nor2 g683(.a(new_n734_), .b(new_n652_), .O(new_n735_));
  inv1 g684(.a(new_n735_), .O(o_5_));
  nor2 g685(.a(new_n441_), .b(new_n432_), .O(new_n737_));
  inv1 g686(.a(new_n737_), .O(new_n738_));
  nor2 g687(.a(new_n738_), .b(new_n420_), .O(new_n739_));
  inv1 g688(.a(new_n739_), .O(new_n740_));
  nor2 g689(.a(new_n740_), .b(new_n532_), .O(new_n741_));
  inv1 g690(.a(new_n741_), .O(new_n742_));
  nor2 g691(.a(new_n647_), .b(new_n413_), .O(new_n743_));
  inv1 g692(.a(new_n743_), .O(new_n744_));
  nor2 g693(.a(new_n744_), .b(new_n742_), .O(new_n745_));
  inv1 g694(.a(new_n745_), .O(o_6_));
  nor2 g695(.a(o_23_), .b(new_n321_), .O(new_n747_));
  inv1 g696(.a(new_n747_), .O(new_n748_));
  nor2 g697(.a(new_n748_), .b(o_13_), .O(new_n749_));
  inv1 g698(.a(new_n749_), .O(new_n750_));
  nor2 g699(.a(new_n750_), .b(new_n723_), .O(new_n751_));
  inv1 g700(.a(new_n751_), .O(o_3_));
  nor2 g701(.a(i_14_), .b(i_20_), .O(o_4_));
endmodule


